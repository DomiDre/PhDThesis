@Filename: C:\vsm-lv\System_Admin\data\Dominique\DD150\empty_sample_holder\empty_sample_holder-Hys-00.VHD
@Measurement Controlfilename: c:\vsm-lv\System_Admin\Recipes\VC_HL_quickscan_allrange.VHC
@Calibration filename: c:\vsm-lv\System_Admin\settings\default.cal
@Parameter Filec:\vsm-lv\System_Admin\settings\default.cal
@Operator: System_Admin
@Samplename: empty_sample_holder
@Date: Friday, October 14, 2016    (2016-10-14)
@Time: 09:32:50
@Test ID: test
@Apparatus: EZ7; LabVSM; Customer: Grubenhagen; first started on: Wednesday February 03, , 2015
[Installed Options]
VSM Model="EV X"
VSM=TRUE    
Torque=FALSE    
Signal Processor="SRS SR 830"
Torque Signal Processor="NI-6210"
Unipolar=FALSE    
Automation=FALSE    
MR=FALSE    
Torque Signal Inversion=TRUE    
VSM DAQ Card=TRUE    
Time Constant="0.1 s"
DAQ Output=FALSE    

[Signal and Coils]
Signal Connection="A-B"
Vector Coils=FALSE    
Stationary Coils=FALSE    
Z Coils=FALSE    
Sensor Angle="0 deg"
Time Between Averages=0.150000    
Y Averages Multiplier=1    
Reference Source="External"
SR830 Frequency=75.000000    

[Rotation]
Automatic Rotation=TRUE    
Rotate Option="Mdrive"
Rotation Display=FALSE    
Max Angle=400.000000    
Min Angle=-400.000000    
Rotation Serial Port=1    
Rotation Display Serial Port=1    
Torque Rotation Serial Port=4    

[Field]
Gaussmeter="32 KP DRC"
Gauss Probe="1 x"
Maximum Field=19000.000000    
Wait Time=4.000000    
Sweeprate Array="1500.000, 500.000, 100.000, 10.000, "
Averaging Array="1, 1, 1, 10, "
Precision Array="3.000, 0.500, 0.200, 0.200, "
Stability Array="1.000, 1.000, 0.500, 0.100, "
FCM-10 Address="GPIB0::16::INSTR"
Minimum Sweep Time=2.000000    
Minimum Sweep Rate Divider=40.000000    
Stability Time Between Readings=0.300000    
Number of Readings for Stability Check=2.000000    
Slow Approach=TRUE    
Slow Start %=90.000000    
Slow Approach Max Sweep Rate Divider=10.000000    
Max Slow Sweep Time=4.000000    

[MR]
MR Signal Processor=Manual VSM
Punch Through="Variable 0-10V"
Automation Comm Port=0
Max Current=20.000000    
Min AD Voltage=4.600000    
Max AD Voltage=7.000000    
MR Option=FALSE    
MS MR Signal Processor=FALSE    
AC&DC Current Source=FALSE    

[Temperature Control]
Temperature Control=TRUE    
Boil Off Nitrogen=FALSE    
Liquid Helium=FALSE    
Leave Temperature On=TRUE    
Temperature Control Type="SI 9700"
Sensor A="E-type"
Sensor B="E-type"
Control Sensor="A"
Sensor A Table=""
Sensor B Table=""
ITC Serial Port=2    
TC GPIB Address=15    
Temperature Log File="/c/vsm-lv/temperature.log"
Default Temperature=298.150000    
Gas Switching Temperature=333.150000    
Default Soak Time=120.000000    
Set Temperature Sample Time=10.000000    
Temperature Accuracy=1.000000    
Temperature Accuracy %=1.000000    
Automatic Gas Switching=FALSE    
1000 C Option=FALSE    
Number of points for accuracy wait=90    
Time between points for accuracy wait=1.000000    
Wait for Heat Exchanger Removal=FALSE    
Removal Temperature=0.000000    
Wait Time for Heat Exchanger Removal=0.000000    

[SI 9700]
P=1    
I=20    
D=0    
HE-P=1    
HE-I=20    
HE-D=0    
Max T Sweep Seed=1.000000
Min T Sweep Seed=0.200000
Max Heater Power=80    
Max T Sweep Speed=60.000000    
Min T Sweep Speed=12.000000    

[Other]
Transverse Direction="Absolute"
Default Transverse Direction=90.000000    
Time Dependence Start Field Distance=10.000000    
Minimum Remanence Wait Time=2.000000    
Default AC Demag Max Field=10000.000000    
AC Demag Minimum Field=1.000000    
Max Lockin Phase Error=90    
Mains Frequency=50.000000    
Samples Per Cycle=100    

[Interlock]
Door Lock=FALSE    
Interlock=FALSE    
Light Tower=FALSE    
Interlock Interface Name="Dev3"

[Torque Interface]
Torque Interface Name="Dev2"

[Exit Gas Heater Settings]
EGH PC Control=FALSE    
EGH Serial Port=0    
EGH Voltages=""

[VSM Interface]
VSM Interface Name="Dev1"

[MR Interface]
MR Interface Name="Dev1"

[DAQ Communication]
Protocol="Mx"
Remove Spikes=TRUE    

[Sensor Table]
1st Column=0    
Temperature Unit=0    

[Communication]
LIA 1 Address="GPIB0::8::INSTR"
LIA 2 Address=""
VSM Rotation Address="COM1"
Torque Rotation Address=""
Rotation Display Address=""
SI9700 Address="COM12"
EGH Address=""
Communication Mode="Original"
LIA Baud Rate="19200"
LIA Serial Read Delay=50    

[LIA]
Local=0    
Minimum Sensitivity="5 uV"

[MR External Current Source]
Ext I Src Adddress=""
AC MR Channel=""
DC MR Channel=""
Read Termination Character="CR"
CS Baud Rate="300"
Flow Control="Off"
Which LIA="1"
Input="A"
Ref Slope="Sine"
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 2.686E-2 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: MicroSense EasyVSM Software version EasyVSM 20150305-01
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to -0.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set VSM DAQ AO0 Voltage to 10.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 2:      Set VSM DAQ AO1 Voltage to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Applied Field to 0.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 4:      Set Auto Range Signal to 10.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = No
@Number of sections= 3
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From:  0.0000 [Oe] To: 19000.0000 [Oe] Min Stepsize/Sweeprate = 1000.0000 [Oe] Max Stepsize/Sweeprate = 1000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Measured Signal(s) = X
@Section 0 END
@Section 1: Hysteresis
@Preparation Actions: None
@Main Parameter Setup:
     From: 19000.0000 [Oe] To: -19000.0000 [Oe] Min Stepsize/Sweeprate = 1000.0000 [Oe] Max Stepsize/Sweeprate = 1000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: -19000.0000 [Oe] To: 19000.0000 [Oe] Min Stepsize/Sweeprate = 1000.0000 [Oe] Max Stepsize/Sweeprate = 1000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 2 END
@@Plot Settings
Number of plots: 1
Plot 0: Hysteresis = On; Section: 0; Signal: X; Label: Hys X; Point style: 2; Interpolation: On; Color: 14417948; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = FALSE
Sensor Angle = 0 deg
@Gauss Range: 30 kOe
@Emu Range: 5 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 5
@Rot 0 deg cal: -21170
@Rot 360 deg cal: 20810
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 10530
@Emu/v: 58.557
@Y Coils Correction Factor: 1.385
@Sample Shape Correction Factor: 1.000
@Coil Angle Alpha: 45.000
@Coil Angle Beta: -45.000
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 17
14997.000000   1.000000
15246.000000   1.000145
15496.000000   1.000446
15746.000000   1.000592
15995.000000   1.000892
16246.000000   1.001261
16495.000000   1.001631
16745.000000   1.002000
16995.000000   1.002448
17245.000000   1.002965
17495.000000   1.003491
17745.000000   1.004009
17994.000000   1.004605
18244.000000   1.005202
18494.000000   1.006025
18744.000000   1.006702
18994.000000   1.007597
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 0.700000
Background Subtraction = Yes   Method = Straight Line
Background slope x, y, z [emu/Oe] = -1.237658E-7   -0.000000E+0   -0.000000E+0
Background Offset x, y, z [emu] = 9.062174E-7   -0.000000E+0   -0.000000E+0
Angular Sensitivity Correction = Yes
Angular Sensitivity array length = 361
0.000000   1.000026E+0   0.000000E+0   0.000000
1.000000   9.998824E-1   0.000000E+0   0.000000
2.000000   9.997501E-1   0.000000E+0   0.000000
3.000000   9.996408E-1   0.000000E+0   0.000000
4.000000   9.995661E-1   0.000000E+0   0.000000
5.000000   9.995373E-1   0.000000E+0   0.000000
6.000000   9.995662E-1   0.000000E+0   0.000000
7.000000   9.996640E-1   0.000000E+0   0.000000
8.000000   9.998424E-1   0.000000E+0   0.000000
9.000000   1.000113E+0   0.000000E+0   0.000000
10.000000   1.000487E+0   0.000000E+0   0.000000
11.000000   1.000976E+0   0.000000E+0   0.000000
12.000000   1.001591E+0   0.000000E+0   0.000000
13.000000   1.002345E+0   0.000000E+0   0.000000
14.000000   1.003248E+0   0.000000E+0   0.000000
15.000000   1.004313E+0   0.000000E+0   0.000000
16.000000   1.005547E+0   0.000000E+0   0.000000
17.000000   1.006952E+0   0.000000E+0   0.000000
18.000000   1.008524E+0   0.000000E+0   0.000000
19.000000   1.010260E+0   0.000000E+0   0.000000
20.000000   1.012158E+0   0.000000E+0   0.000000
21.000000   1.014215E+0   0.000000E+0   0.000000
22.000000   1.016429E+0   0.000000E+0   0.000000
23.000000   1.018797E+0   0.000000E+0   0.000000
24.000000   1.021316E+0   0.000000E+0   0.000000
25.000000   1.023983E+0   0.000000E+0   0.000000
26.000000   1.026796E+0   0.000000E+0   0.000000
27.000000   1.029751E+0   0.000000E+0   0.000000
28.000000   1.032848E+0   0.000000E+0   0.000000
29.000000   1.036082E+0   0.000000E+0   0.000000
30.000000   1.039451E+0   0.000000E+0   0.000000
31.000000   1.042951E+0   0.000000E+0   0.000000
32.000000   1.046574E+0   0.000000E+0   0.000000
33.000000   1.050309E+0   0.000000E+0   0.000000
34.000000   1.054148E+0   0.000000E+0   0.000000
35.000000   1.058079E+0   0.000000E+0   0.000000
36.000000   1.062094E+0   0.000000E+0   0.000000
37.000000   1.066183E+0   0.000000E+0   0.000000
38.000000   1.070335E+0   0.000000E+0   0.000000
39.000000   1.074542E+0   0.000000E+0   0.000000
40.000000   1.078793E+0   0.000000E+0   0.000000
41.000000   1.083078E+0   0.000000E+0   0.000000
42.000000   1.087388E+0   0.000000E+0   0.000000
43.000000   1.091713E+0   0.000000E+0   0.000000
44.000000   1.096043E+0   0.000000E+0   0.000000
45.000000   1.100369E+0   0.000000E+0   0.000000
46.000000   1.104681E+0   0.000000E+0   0.000000
47.000000   1.108977E+0   0.000000E+0   0.000000
48.000000   1.113255E+0   0.000000E+0   0.000000
49.000000   1.117512E+0   0.000000E+0   0.000000
50.000000   1.121748E+0   0.000000E+0   0.000000
51.000000   1.125960E+0   0.000000E+0   0.000000
52.000000   1.130146E+0   0.000000E+0   0.000000
53.000000   1.134304E+0   0.000000E+0   0.000000
54.000000   1.138432E+0   0.000000E+0   0.000000
55.000000   1.142529E+0   0.000000E+0   0.000000
56.000000   1.146593E+0   0.000000E+0   0.000000
57.000000   1.150621E+0   0.000000E+0   0.000000
58.000000   1.154612E+0   0.000000E+0   0.000000
59.000000   1.158564E+0   0.000000E+0   0.000000
60.000000   1.162475E+0   0.000000E+0   0.000000
61.000000   1.166339E+0   0.000000E+0   0.000000
62.000000   1.170133E+0   0.000000E+0   0.000000
63.000000   1.173831E+0   0.000000E+0   0.000000
64.000000   1.177406E+0   0.000000E+0   0.000000
65.000000   1.180831E+0   0.000000E+0   0.000000
66.000000   1.184079E+0   0.000000E+0   0.000000
67.000000   1.187125E+0   0.000000E+0   0.000000
68.000000   1.189940E+0   0.000000E+0   0.000000
69.000000   1.192499E+0   0.000000E+0   0.000000
70.000000   1.194775E+0   0.000000E+0   0.000000
71.000000   1.196740E+0   0.000000E+0   0.000000
72.000000   1.198369E+0   0.000000E+0   0.000000
73.000000   1.199634E+0   0.000000E+0   0.000000
74.000000   1.200509E+0   0.000000E+0   0.000000
75.000000   1.200967E+0   0.000000E+0   0.000000
76.000000   1.200994E+0   0.000000E+0   0.000000
77.000000   1.200624E+0   0.000000E+0   0.000000
78.000000   1.199905E+0   0.000000E+0   0.000000
79.000000   1.198883E+0   0.000000E+0   0.000000
80.000000   1.197605E+0   0.000000E+0   0.000000
81.000000   1.196119E+0   0.000000E+0   0.000000
82.000000   1.194472E+0   0.000000E+0   0.000000
83.000000   1.192710E+0   0.000000E+0   0.000000
84.000000   1.190880E+0   0.000000E+0   0.000000
85.000000   1.189031E+0   0.000000E+0   0.000000
86.000000   1.187207E+0   0.000000E+0   0.000000
87.000000   1.185457E+0   0.000000E+0   0.000000
88.000000   1.183828E+0   0.000000E+0   0.000000
89.000000   1.182367E+0   0.000000E+0   0.000000
90.000000   1.181120E+0   0.000000E+0   0.000000
91.000000   1.180125E+0   0.000000E+0   0.000000
92.000000   1.179386E+0   0.000000E+0   0.000000
93.000000   1.178896E+0   0.000000E+0   0.000000
94.000000   1.178648E+0   0.000000E+0   0.000000
95.000000   1.178636E+0   0.000000E+0   0.000000
96.000000   1.178854E+0   0.000000E+0   0.000000
97.000000   1.179294E+0   0.000000E+0   0.000000
98.000000   1.179952E+0   0.000000E+0   0.000000
99.000000   1.180819E+0   0.000000E+0   0.000000
100.000000   1.181891E+0   0.000000E+0   0.000000
101.000000   1.183160E+0   0.000000E+0   0.000000
102.000000   1.184620E+0   0.000000E+0   0.000000
103.000000   1.186264E+0   0.000000E+0   0.000000
104.000000   1.188087E+0   0.000000E+0   0.000000
105.000000   1.190081E+0   0.000000E+0   0.000000
106.000000   1.192236E+0   0.000000E+0   0.000000
107.000000   1.194518E+0   0.000000E+0   0.000000
108.000000   1.196891E+0   0.000000E+0   0.000000
109.000000   1.199318E+0   0.000000E+0   0.000000
110.000000   1.201761E+0   0.000000E+0   0.000000
111.000000   1.204182E+0   0.000000E+0   0.000000
112.000000   1.206545E+0   0.000000E+0   0.000000
113.000000   1.208812E+0   0.000000E+0   0.000000
114.000000   1.210946E+0   0.000000E+0   0.000000
115.000000   1.212909E+0   0.000000E+0   0.000000
116.000000   1.214664E+0   0.000000E+0   0.000000
117.000000   1.216174E+0   0.000000E+0   0.000000
118.000000   1.217402E+0   0.000000E+0   0.000000
119.000000   1.218310E+0   0.000000E+0   0.000000
120.000000   1.218860E+0   0.000000E+0   0.000000
121.000000   1.219027E+0   0.000000E+0   0.000000
122.000000   1.218821E+0   0.000000E+0   0.000000
123.000000   1.218265E+0   0.000000E+0   0.000000
124.000000   1.217382E+0   0.000000E+0   0.000000
125.000000   1.216194E+0   0.000000E+0   0.000000
126.000000   1.214723E+0   0.000000E+0   0.000000
127.000000   1.212992E+0   0.000000E+0   0.000000
128.000000   1.211022E+0   0.000000E+0   0.000000
129.000000   1.208837E+0   0.000000E+0   0.000000
130.000000   1.206459E+0   0.000000E+0   0.000000
131.000000   1.203910E+0   0.000000E+0   0.000000
132.000000   1.201212E+0   0.000000E+0   0.000000
133.000000   1.198388E+0   0.000000E+0   0.000000
134.000000   1.195459E+0   0.000000E+0   0.000000
135.000000   1.192449E+0   0.000000E+0   0.000000
136.000000   1.189376E+0   0.000000E+0   0.000000
137.000000   1.186243E+0   0.000000E+0   0.000000
138.000000   1.183050E+0   0.000000E+0   0.000000
139.000000   1.179797E+0   0.000000E+0   0.000000
140.000000   1.176482E+0   0.000000E+0   0.000000
141.000000   1.173105E+0   0.000000E+0   0.000000
142.000000   1.169667E+0   0.000000E+0   0.000000
143.000000   1.166166E+0   0.000000E+0   0.000000
144.000000   1.162602E+0   0.000000E+0   0.000000
145.000000   1.158975E+0   0.000000E+0   0.000000
146.000000   1.155283E+0   0.000000E+0   0.000000
147.000000   1.151528E+0   0.000000E+0   0.000000
148.000000   1.147707E+0   0.000000E+0   0.000000
149.000000   1.143822E+0   0.000000E+0   0.000000
150.000000   1.139870E+0   0.000000E+0   0.000000
151.000000   1.135854E+0   0.000000E+0   0.000000
152.000000   1.131784E+0   0.000000E+0   0.000000
153.000000   1.127671E+0   0.000000E+0   0.000000
154.000000   1.123527E+0   0.000000E+0   0.000000
155.000000   1.119362E+0   0.000000E+0   0.000000
156.000000   1.115190E+0   0.000000E+0   0.000000
157.000000   1.111022E+0   0.000000E+0   0.000000
158.000000   1.106868E+0   0.000000E+0   0.000000
159.000000   1.102742E+0   0.000000E+0   0.000000
160.000000   1.098653E+0   0.000000E+0   0.000000
161.000000   1.094615E+0   0.000000E+0   0.000000
162.000000   1.090639E+0   0.000000E+0   0.000000
163.000000   1.086736E+0   0.000000E+0   0.000000
164.000000   1.082918E+0   0.000000E+0   0.000000
165.000000   1.079196E+0   0.000000E+0   0.000000
166.000000   1.075581E+0   0.000000E+0   0.000000
167.000000   1.072078E+0   0.000000E+0   0.000000
168.000000   1.068691E+0   0.000000E+0   0.000000
169.000000   1.065422E+0   0.000000E+0   0.000000
170.000000   1.062276E+0   0.000000E+0   0.000000
171.000000   1.059256E+0   0.000000E+0   0.000000
172.000000   1.056366E+0   0.000000E+0   0.000000
173.000000   1.053609E+0   0.000000E+0   0.000000
174.000000   1.050989E+0   0.000000E+0   0.000000
175.000000   1.048510E+0   0.000000E+0   0.000000
176.000000   1.046174E+0   0.000000E+0   0.000000
177.000000   1.043987E+0   0.000000E+0   0.000000
178.000000   1.041950E+0   0.000000E+0   0.000000
179.000000   1.040068E+0   0.000000E+0   0.000000
180.000000   1.038345E+0   0.000000E+0   0.000000
181.000000   1.036783E+0   0.000000E+0   0.000000
182.000000   1.035385E+0   0.000000E+0   0.000000
183.000000   1.034152E+0   0.000000E+0   0.000000
184.000000   1.033086E+0   0.000000E+0   0.000000
185.000000   1.032187E+0   0.000000E+0   0.000000
186.000000   1.031459E+0   0.000000E+0   0.000000
187.000000   1.030901E+0   0.000000E+0   0.000000
188.000000   1.030516E+0   0.000000E+0   0.000000
189.000000   1.030306E+0   0.000000E+0   0.000000
190.000000   1.030271E+0   0.000000E+0   0.000000
191.000000   1.030414E+0   0.000000E+0   0.000000
192.000000   1.030736E+0   0.000000E+0   0.000000
193.000000   1.031238E+0   0.000000E+0   0.000000
194.000000   1.031922E+0   0.000000E+0   0.000000
195.000000   1.032790E+0   0.000000E+0   0.000000
196.000000   1.033841E+0   0.000000E+0   0.000000
197.000000   1.035069E+0   0.000000E+0   0.000000
198.000000   1.036465E+0   0.000000E+0   0.000000
199.000000   1.038023E+0   0.000000E+0   0.000000
200.000000   1.039733E+0   0.000000E+0   0.000000
201.000000   1.041588E+0   0.000000E+0   0.000000
202.000000   1.043579E+0   0.000000E+0   0.000000
203.000000   1.045699E+0   0.000000E+0   0.000000
204.000000   1.047938E+0   0.000000E+0   0.000000
205.000000   1.050290E+0   0.000000E+0   0.000000
206.000000   1.052746E+0   0.000000E+0   0.000000
207.000000   1.055298E+0   0.000000E+0   0.000000
208.000000   1.057938E+0   0.000000E+0   0.000000
209.000000   1.060657E+0   0.000000E+0   0.000000
210.000000   1.063448E+0   0.000000E+0   0.000000
211.000000   1.066303E+0   0.000000E+0   0.000000
212.000000   1.069213E+0   0.000000E+0   0.000000
213.000000   1.072170E+0   0.000000E+0   0.000000
214.000000   1.075167E+0   0.000000E+0   0.000000
215.000000   1.078196E+0   0.000000E+0   0.000000
216.000000   1.081247E+0   0.000000E+0   0.000000
217.000000   1.084314E+0   0.000000E+0   0.000000
218.000000   1.087389E+0   0.000000E+0   0.000000
219.000000   1.090463E+0   0.000000E+0   0.000000
220.000000   1.093528E+0   0.000000E+0   0.000000
221.000000   1.096576E+0   0.000000E+0   0.000000
222.000000   1.099599E+0   0.000000E+0   0.000000
223.000000   1.102590E+0   0.000000E+0   0.000000
224.000000   1.105540E+0   0.000000E+0   0.000000
225.000000   1.108441E+0   0.000000E+0   0.000000
226.000000   1.111288E+0   0.000000E+0   0.000000
227.000000   1.114083E+0   0.000000E+0   0.000000
228.000000   1.116834E+0   0.000000E+0   0.000000
229.000000   1.119546E+0   0.000000E+0   0.000000
230.000000   1.122224E+0   0.000000E+0   0.000000
231.000000   1.124876E+0   0.000000E+0   0.000000
232.000000   1.127507E+0   0.000000E+0   0.000000
233.000000   1.130123E+0   0.000000E+0   0.000000
234.000000   1.132730E+0   0.000000E+0   0.000000
235.000000   1.135334E+0   0.000000E+0   0.000000
236.000000   1.137940E+0   0.000000E+0   0.000000
237.000000   1.140556E+0   0.000000E+0   0.000000
238.000000   1.143186E+0   0.000000E+0   0.000000
239.000000   1.145838E+0   0.000000E+0   0.000000
240.000000   1.148516E+0   0.000000E+0   0.000000
241.000000   1.151221E+0   0.000000E+0   0.000000
242.000000   1.153928E+0   0.000000E+0   0.000000
243.000000   1.156608E+0   0.000000E+0   0.000000
244.000000   1.159229E+0   0.000000E+0   0.000000
245.000000   1.161761E+0   0.000000E+0   0.000000
246.000000   1.164173E+0   0.000000E+0   0.000000
247.000000   1.166436E+0   0.000000E+0   0.000000
248.000000   1.168519E+0   0.000000E+0   0.000000
249.000000   1.170391E+0   0.000000E+0   0.000000
250.000000   1.172022E+0   0.000000E+0   0.000000
251.000000   1.173381E+0   0.000000E+0   0.000000
252.000000   1.174439E+0   0.000000E+0   0.000000
253.000000   1.175164E+0   0.000000E+0   0.000000
254.000000   1.175526E+0   0.000000E+0   0.000000
255.000000   1.175494E+0   0.000000E+0   0.000000
256.000000   1.175054E+0   0.000000E+0   0.000000
257.000000   1.174243E+0   0.000000E+0   0.000000
258.000000   1.173118E+0   0.000000E+0   0.000000
259.000000   1.171731E+0   0.000000E+0   0.000000
260.000000   1.170138E+0   0.000000E+0   0.000000
261.000000   1.168393E+0   0.000000E+0   0.000000
262.000000   1.166549E+0   0.000000E+0   0.000000
263.000000   1.164661E+0   0.000000E+0   0.000000
264.000000   1.162784E+0   0.000000E+0   0.000000
265.000000   1.160972E+0   0.000000E+0   0.000000
266.000000   1.159278E+0   0.000000E+0   0.000000
267.000000   1.157758E+0   0.000000E+0   0.000000
268.000000   1.156464E+0   0.000000E+0   0.000000
269.000000   1.155453E+0   0.000000E+0   0.000000
270.000000   1.154778E+0   0.000000E+0   0.000000
271.000000   1.154479E+0   0.000000E+0   0.000000
272.000000   1.154546E+0   0.000000E+0   0.000000
273.000000   1.154954E+0   0.000000E+0   0.000000
274.000000   1.155676E+0   0.000000E+0   0.000000
275.000000   1.156690E+0   0.000000E+0   0.000000
276.000000   1.157968E+0   0.000000E+0   0.000000
277.000000   1.159488E+0   0.000000E+0   0.000000
278.000000   1.161223E+0   0.000000E+0   0.000000
279.000000   1.163148E+0   0.000000E+0   0.000000
280.000000   1.165240E+0   0.000000E+0   0.000000
281.000000   1.167472E+0   0.000000E+0   0.000000
282.000000   1.169820E+0   0.000000E+0   0.000000
283.000000   1.172260E+0   0.000000E+0   0.000000
284.000000   1.174765E+0   0.000000E+0   0.000000
285.000000   1.177311E+0   0.000000E+0   0.000000
286.000000   1.179873E+0   0.000000E+0   0.000000
287.000000   1.182423E+0   0.000000E+0   0.000000
288.000000   1.184933E+0   0.000000E+0   0.000000
289.000000   1.187376E+0   0.000000E+0   0.000000
290.000000   1.189723E+0   0.000000E+0   0.000000
291.000000   1.191947E+0   0.000000E+0   0.000000
292.000000   1.194019E+0   0.000000E+0   0.000000
293.000000   1.195912E+0   0.000000E+0   0.000000
294.000000   1.197597E+0   0.000000E+0   0.000000
295.000000   1.199047E+0   0.000000E+0   0.000000
296.000000   1.200234E+0   0.000000E+0   0.000000
297.000000   1.201130E+0   0.000000E+0   0.000000
298.000000   1.201706E+0   0.000000E+0   0.000000
299.000000   1.201936E+0   0.000000E+0   0.000000
300.000000   1.201791E+0   0.000000E+0   0.000000
301.000000   1.201251E+0   0.000000E+0   0.000000
302.000000   1.200329E+0   0.000000E+0   0.000000
303.000000   1.199047E+0   0.000000E+0   0.000000
304.000000   1.197426E+0   0.000000E+0   0.000000
305.000000   1.195488E+0   0.000000E+0   0.000000
306.000000   1.193253E+0   0.000000E+0   0.000000
307.000000   1.190744E+0   0.000000E+0   0.000000
308.000000   1.187980E+0   0.000000E+0   0.000000
309.000000   1.184985E+0   0.000000E+0   0.000000
310.000000   1.181778E+0   0.000000E+0   0.000000
311.000000   1.178381E+0   0.000000E+0   0.000000
312.000000   1.174816E+0   0.000000E+0   0.000000
313.000000   1.171104E+0   0.000000E+0   0.000000
314.000000   1.167266E+0   0.000000E+0   0.000000
315.000000   1.163324E+0   0.000000E+0   0.000000
316.000000   1.159296E+0   0.000000E+0   0.000000
317.000000   1.155191E+0   0.000000E+0   0.000000
318.000000   1.151016E+0   0.000000E+0   0.000000
319.000000   1.146778E+0   0.000000E+0   0.000000
320.000000   1.142484E+0   0.000000E+0   0.000000
321.000000   1.138139E+0   0.000000E+0   0.000000
322.000000   1.133751E+0   0.000000E+0   0.000000
323.000000   1.129325E+0   0.000000E+0   0.000000
324.000000   1.124870E+0   0.000000E+0   0.000000
325.000000   1.120390E+0   0.000000E+0   0.000000
326.000000   1.115894E+0   0.000000E+0   0.000000
327.000000   1.111387E+0   0.000000E+0   0.000000
328.000000   1.106877E+0   0.000000E+0   0.000000
329.000000   1.102369E+0   0.000000E+0   0.000000
330.000000   1.097870E+0   0.000000E+0   0.000000
331.000000   1.093388E+0   0.000000E+0   0.000000
332.000000   1.088932E+0   0.000000E+0   0.000000
333.000000   1.084513E+0   0.000000E+0   0.000000
334.000000   1.080140E+0   0.000000E+0   0.000000
335.000000   1.075824E+0   0.000000E+0   0.000000
336.000000   1.071575E+0   0.000000E+0   0.000000
337.000000   1.067403E+0   0.000000E+0   0.000000
338.000000   1.063319E+0   0.000000E+0   0.000000
339.000000   1.059332E+0   0.000000E+0   0.000000
340.000000   1.055454E+0   0.000000E+0   0.000000
341.000000   1.051693E+0   0.000000E+0   0.000000
342.000000   1.048060E+0   0.000000E+0   0.000000
343.000000   1.044566E+0   0.000000E+0   0.000000
344.000000   1.041221E+0   0.000000E+0   0.000000
345.000000   1.038035E+0   0.000000E+0   0.000000
346.000000   1.035014E+0   0.000000E+0   0.000000
347.000000   1.032151E+0   0.000000E+0   0.000000
348.000000   1.029434E+0   0.000000E+0   0.000000
349.000000   1.026853E+0   0.000000E+0   0.000000
350.000000   1.024396E+0   0.000000E+0   0.000000
351.000000   1.022052E+0   0.000000E+0   0.000000
352.000000   1.019809E+0   0.000000E+0   0.000000
353.000000   1.017656E+0   0.000000E+0   0.000000
354.000000   1.015583E+0   0.000000E+0   0.000000
355.000000   1.013576E+0   0.000000E+0   0.000000
356.000000   1.011627E+0   0.000000E+0   0.000000
357.000000   1.009722E+0   0.000000E+0   0.000000
358.000000   1.007851E+0   0.000000E+0   0.000000
359.000000   1.006003E+0   0.000000E+0   0.000000
360.000000   1.004166E+0   0.000000E+0   0.000000
Remove Slope = No

Remove Signal Offset = No
Remove Signal Drift = FALSE; Drift # Points = 0
Remove Field Offset = No
Field Offset Method = Automatic
Field Offset = 0.0000
Remove Field Lag = No
Field Lag Method = Automatic
Field Lag = 0.0000
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0   Filter Type = Median
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = Tuesday, October 11, 2016  10:51:58
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 3
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Temperature 2, Sample Temperature [degC]
Column 4: Raw Applied Field, Applied Field [Oe]
Column 5: Applied Field, Applied Field [Oe]
Column 6: Field Angle, Field Angle [deg]
Column 7: Raw Applied Field For Plot , Applied Field [Oe]
Column 8: Applied Field For Plot , Applied Field [Oe]
Column 9: Raw Signal Mx, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Temperature_2   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Signal_X_direction      
@Time at start of measurement: 09:32:51
@@Data
New Section: Section 0: 
3.541000E+0   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   6.789638E-4   -2.272359E-7   
1.263300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.960000E+2   9.960000E+2   -1.308987E-1   -8.537596E-6   
2.187700E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.997000E+3   1.997000E+3   -2.633190E-1   -1.707172E-5   
3.204200E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.997000E+3   2.997000E+3   -4.020888E-1   -3.207942E-5   
4.129000E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.998000E+3   3.998000E+3   -5.276030E-1   -3.370731E-5   
5.196000E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.998000E+3   4.998000E+3   -6.579794E-1   -4.032129E-5   
6.121400E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.998000E+3   5.998000E+3   -7.890502E-1   -4.762965E-5   
7.094100E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.998000E+3   6.998000E+3   -9.266020E-1   -6.141922E-5   
8.013100E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.998000E+3   7.998000E+3   -1.051684E+0   -6.273826E-5   
9.079300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.998000E+3   8.998000E+3   -1.185862E+0   -7.315488E-5   
9.980300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.998000E+3   9.998000E+3   -1.312426E+0   -7.595543E-5   
1.093890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.099800E+4   1.099800E+4   -1.445863E+0   -8.563071E-5   
1.192530E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.199800E+4   1.199800E+4   -1.567825E+0   -8.382977E-5   
1.291170E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.299800E+4   1.299800E+4   -1.701000E+0   -9.324271E-5   
1.389770E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.399800E+4   1.399800E+4   -1.825325E+0   -9.380517E-5   
1.493350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499800E+4   1.499800E+4   -1.954791E+0   -9.951050E-5   
1.599000E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.599800E+4   1.599800E+4   -2.071408E+0   -9.475178E-5   
1.712640E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.699800E+4   1.699800E+4   -2.201442E+0   -1.055829E-4   
1.826220E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.799700E+4   1.799700E+4   -2.316664E+0   -1.039705E-4   
1.944950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.899600E+4   1.899600E+4   -2.428330E+0   -1.020111E-4   
2.076600E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.800300E+4   1.800300E+4   -2.316357E+0   -1.029633E-4   
2.189730E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700300E+4   1.700300E+4   -2.203320E+0   -1.068757E-4   
2.292920E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600500E+4   1.600500E+4   -2.074506E+0   -9.701361E-5   
2.396650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.500300E+4   1.500300E+4   -1.947221E+0   -9.132856E-5   
2.499890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400300E+4   1.400300E+4   -1.827724E+0   -9.558488E-5   
2.603050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300200E+4   1.300200E+4   -1.701654E+0   -9.340115E-5   
2.701310E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200200E+4   1.200200E+4   -1.575023E+0   -9.053267E-5   
2.799730E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100100E+4   1.100100E+4   -1.449180E+0   -8.857615E-5   
2.897830E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000200E+4   1.000200E+4   -1.312011E+0   -7.504578E-5   
2.991450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.002000E+3   9.002000E+3   -1.185250E+0   -7.204730E-5   
3.088310E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.002000E+3   8.002000E+3   -1.052382E+0   -6.294121E-5   
3.182340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.001000E+3   7.001000E+3   -9.274077E-1   -6.185368E-5   
3.273890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.002000E+3   6.002000E+3   -7.944924E-1   -5.257698E-5   
3.368020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.001000E+3   5.001000E+3   -6.640447E-1   -4.601544E-5   
3.460370E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.002000E+3   4.002000E+3   -5.278158E-1   -3.342505E-5   
3.550140E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.002000E+3   3.002000E+3   -3.965589E-1   -2.593048E-5   
3.642460E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.002000E+3   2.002000E+3   -2.612247E-1   -1.435862E-5   
3.731880E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.001000E+3   1.001000E+3   -1.319539E-1   -8.973984E-6   
3.818940E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.000000E+0   2.000000E+0   -2.225043E-3   -2.883787E-6   
3.909960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.970000E+2   -9.970000E+2   1.292708E-1   4.973479E-6   
4.002530E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.997000E+3   -1.997000E+3   2.639733E-1   1.591361E-5   
4.099440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.998000E+3   -2.998000E+3   3.967117E-1   2.476594E-5   
4.191440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.997000E+3   -3.997000E+3   5.294736E-1   3.388923E-5   
4.285500E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.998000E+3   -4.998000E+3   6.580883E-1   3.861777E-5   
4.382420E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.998000E+3   -5.998000E+3   7.903033E-1   4.707036E-5   
4.476440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.998000E+3   -6.998000E+3   9.211492E-1   5.415385E-5   
4.573280E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.998000E+3   -7.998000E+3   1.043176E+0   5.241850E-5   
4.670220E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.998000E+3   -8.998000E+3   1.182720E+0   6.820022E-5   
4.764210E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.998000E+3   -9.998000E+3   1.303984E+0   6.570126E-5   
4.859790E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.099800E+4   -1.099800E+4   1.439123E+0   7.707824E-5   
4.958550E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.199800E+4   -1.199800E+4   1.569069E+0   8.326111E-5   
5.054390E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.299900E+4   -1.299900E+4   1.698600E+0   8.890680E-5   
5.153140E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.399700E+4   -1.399700E+4   1.820895E+0   8.768599E-5   
5.256990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.499800E+4   -1.499800E+4   1.950755E+0   9.366107E-5   
5.365850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.599800E+4   -1.599800E+4   2.069685E+0   9.121502E-5   
5.474810E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.699800E+4   -1.699800E+4   2.196753E+0   9.906957E-5   
5.588630E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.799700E+4   -1.799700E+4   2.311189E+0   9.665762E-5   
5.717680E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.899900E+4   -1.899900E+4   2.425188E+0   9.666211E-5   
5.844650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.800400E+4   -1.800400E+4   2.312432E+0   9.709052E-5   
5.958120E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.700400E+4   -1.700400E+4   2.199566E+0   1.011826E-4   
6.066570E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.600300E+4   -1.600300E+4   2.078194E+0   9.913212E-5   
6.169960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.500300E+4   -1.500300E+4   1.949992E+0   9.228711E-5   
6.273430E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.400200E+4   -1.400200E+4   1.825085E+0   9.125759E-5   
6.376880E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.300300E+4   -1.300300E+4   1.694521E+0   8.433257E-5   
6.475370E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.200200E+4   -1.200200E+4   1.571599E+0   8.529693E-5   
6.573930E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.100200E+4   -1.100200E+4   1.439406E+0   7.686543E-5   
6.667270E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000100E+4   -1.000100E+4   1.311947E+0   7.329270E-5   
6.760950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.002000E+3   -9.002000E+3   1.186908E+0   7.189323E-5   
6.857550E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.001000E+3   -8.001000E+3   1.056461E+0   6.533169E-5   
6.954170E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.002000E+3   -7.002000E+3   9.217582E-1   5.426780E-5   
7.043090E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.002000E+3   -6.002000E+3   7.937722E-1   5.004428E-5   
7.139850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.001000E+3   -5.001000E+3   6.605758E-1   4.073403E-5   
7.231780E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.001000E+3   -4.001000E+3   5.298007E-1   3.372127E-5   
7.320730E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.002000E+3   -3.002000E+3   3.962100E-1   2.376915E-5   
7.412590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.001000E+3   -2.001000E+3   2.656530E-1   1.709835E-5   
7.504580E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.002000E+3   -1.002000E+3   1.298161E-1   4.899944E-6   
7.591140E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.000000E+0   -2.000000E+0   2.617691E-4   -8.919731E-7   
7.682030E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.960000E+2   9.960000E+2   -1.309068E-1   -8.545677E-6   
7.774490E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.998000E+3   1.998000E+3   -2.633843E-1   -1.701330E-5   
7.866860E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.997000E+3   2.997000E+3   -3.982823E-1   -2.827279E-5   
7.959290E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.998000E+3   3.998000E+3   -5.318295E-1   -3.793392E-5   
8.056660E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.998000E+3   4.998000E+3   -6.597045E-1   -4.204641E-5   
8.153990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.998000E+3   5.998000E+3   -7.862465E-1   -4.482589E-5   
8.251330E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.998000E+3   6.998000E+3   -9.171345E-1   -5.195154E-5   
8.343200E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.999000E+3   7.999000E+3   -1.055566E+0   -6.649689E-5   
8.440510E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.998000E+3   8.998000E+3   -1.171420E+0   -5.871210E-5   
8.532380E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.998000E+3   9.998000E+3   -1.312121E+0   -7.565093E-5   
8.627710E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.099800E+4   1.099800E+4   -1.443616E+0   -8.338325E-5   
8.726350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.199900E+4   1.199900E+4   -1.572123E+0   -8.800417E-5   
8.824990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.299800E+4   1.299800E+4   -1.699580E+0   -9.182209E-5   
8.923640E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.399800E+4   1.399800E+4   -1.823908E+0   -9.238806E-5   
9.027320E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499800E+4   1.499800E+4   -1.951977E+0   -9.669620E-5   
9.132910E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.599900E+4   1.599900E+4   -2.068005E+0   -9.122551E-5   
9.246550E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.699800E+4   1.699800E+4   -2.196467E+0   -1.005955E-4   
9.360250E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.799700E+4   1.799700E+4   -2.309749E+0   -9.702289E-5   
9.483960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.899700E+4   1.899700E+4   -2.428571E+0   -1.021295E-4   
@@END Data.
@Time at end of measurement: 09:48:42
@Instrument  Changes:
@Emu Range: 50 uV
@END Instrument  Changes:
@@Final Manipulated Data
New Section: Section 0: 
3.541000E+0   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   6.789638E-4   -2.272359E-7   
1.263300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.960000E+2   9.960000E+2   -1.308987E-1   -8.537596E-6   
2.187700E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.997000E+3   1.997000E+3   -2.633190E-1   -1.707172E-5   
3.204200E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.997000E+3   2.997000E+3   -4.020888E-1   -3.207942E-5   
4.129000E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.998000E+3   3.998000E+3   -5.276030E-1   -3.370731E-5   
5.196000E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.998000E+3   4.998000E+3   -6.579794E-1   -4.032129E-5   
6.121400E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.998000E+3   5.998000E+3   -7.890502E-1   -4.762965E-5   
7.094100E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.998000E+3   6.998000E+3   -9.266020E-1   -6.141922E-5   
8.013100E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.998000E+3   7.998000E+3   -1.051684E+0   -6.273826E-5   
9.079300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.998000E+3   8.998000E+3   -1.185862E+0   -7.315488E-5   
9.980300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.998000E+3   9.998000E+3   -1.312426E+0   -7.595543E-5   
1.093890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.099800E+4   1.099800E+4   -1.445863E+0   -8.563071E-5   
1.192530E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.199800E+4   1.199800E+4   -1.567825E+0   -8.382977E-5   
1.291170E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.299800E+4   1.299800E+4   -1.701000E+0   -9.324271E-5   
1.389770E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.399800E+4   1.399800E+4   -1.825325E+0   -9.380517E-5   
1.493350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499800E+4   1.499800E+4   -1.954791E+0   -9.951050E-5   
1.599000E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.599800E+4   1.599800E+4   -2.071408E+0   -9.475178E-5   
1.712640E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.699800E+4   1.699800E+4   -2.201442E+0   -1.055829E-4   
1.826220E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.799700E+4   1.799700E+4   -2.316664E+0   -1.039705E-4   
1.944950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.899600E+4   1.899600E+4   -2.428330E+0   -1.020111E-4   
2.076600E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.800300E+4   1.800300E+4   -2.316357E+0   -1.029633E-4   
2.189730E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700300E+4   1.700300E+4   -2.203320E+0   -1.068757E-4   
2.292920E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600500E+4   1.600500E+4   -2.074506E+0   -9.701361E-5   
2.396650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.500300E+4   1.500300E+4   -1.947221E+0   -9.132856E-5   
2.499890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400300E+4   1.400300E+4   -1.827724E+0   -9.558488E-5   
2.603050E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300200E+4   1.300200E+4   -1.701654E+0   -9.340115E-5   
2.701310E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200200E+4   1.200200E+4   -1.575023E+0   -9.053267E-5   
2.799730E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100100E+4   1.100100E+4   -1.449180E+0   -8.857615E-5   
2.897830E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000200E+4   1.000200E+4   -1.312011E+0   -7.504578E-5   
2.991450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.002000E+3   9.002000E+3   -1.185250E+0   -7.204730E-5   
3.088310E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.002000E+3   8.002000E+3   -1.052382E+0   -6.294121E-5   
3.182340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.001000E+3   7.001000E+3   -9.274077E-1   -6.185368E-5   
3.273890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.002000E+3   6.002000E+3   -7.944924E-1   -5.257698E-5   
3.368020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.001000E+3   5.001000E+3   -6.640447E-1   -4.601544E-5   
3.460370E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.002000E+3   4.002000E+3   -5.278158E-1   -3.342505E-5   
3.550140E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.002000E+3   3.002000E+3   -3.965589E-1   -2.593048E-5   
3.642460E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.002000E+3   2.002000E+3   -2.612247E-1   -1.435862E-5   
3.731880E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.001000E+3   1.001000E+3   -1.319539E-1   -8.973984E-6   
3.818940E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.000000E+0   2.000000E+0   -2.225043E-3   -2.883787E-6   
3.909960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.970000E+2   -9.970000E+2   1.292708E-1   4.973479E-6   
4.002530E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.997000E+3   -1.997000E+3   2.639733E-1   1.591361E-5   
4.099440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.998000E+3   -2.998000E+3   3.967117E-1   2.476594E-5   
4.191440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.997000E+3   -3.997000E+3   5.294736E-1   3.388923E-5   
4.285500E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.998000E+3   -4.998000E+3   6.580883E-1   3.861777E-5   
4.382420E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.998000E+3   -5.998000E+3   7.903033E-1   4.707036E-5   
4.476440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.998000E+3   -6.998000E+3   9.211492E-1   5.415385E-5   
4.573280E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.998000E+3   -7.998000E+3   1.043176E+0   5.241850E-5   
4.670220E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.998000E+3   -8.998000E+3   1.182720E+0   6.820022E-5   
4.764210E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.998000E+3   -9.998000E+3   1.303984E+0   6.570126E-5   
4.859790E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.099800E+4   -1.099800E+4   1.439123E+0   7.707824E-5   
4.958550E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.199800E+4   -1.199800E+4   1.569069E+0   8.326111E-5   
5.054390E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.299900E+4   -1.299900E+4   1.698600E+0   8.890680E-5   
5.153140E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.399700E+4   -1.399700E+4   1.820895E+0   8.768599E-5   
5.256990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.499800E+4   -1.499800E+4   1.950755E+0   9.366107E-5   
5.365850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.599800E+4   -1.599800E+4   2.069685E+0   9.121502E-5   
5.474810E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.699800E+4   -1.699800E+4   2.196753E+0   9.906957E-5   
5.588630E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.799700E+4   -1.799700E+4   2.311189E+0   9.665762E-5   
5.717680E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.899900E+4   -1.899900E+4   2.425188E+0   9.666211E-5   
5.844650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.800400E+4   -1.800400E+4   2.312432E+0   9.709052E-5   
5.958120E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.700400E+4   -1.700400E+4   2.199566E+0   1.011826E-4   
6.066570E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.600300E+4   -1.600300E+4   2.078194E+0   9.913212E-5   
6.169960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.500300E+4   -1.500300E+4   1.949992E+0   9.228711E-5   
6.273430E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.400200E+4   -1.400200E+4   1.825085E+0   9.125759E-5   
6.376880E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.300300E+4   -1.300300E+4   1.694521E+0   8.433257E-5   
6.475370E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.200200E+4   -1.200200E+4   1.571599E+0   8.529693E-5   
6.573930E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.100200E+4   -1.100200E+4   1.439406E+0   7.686543E-5   
6.667270E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000100E+4   -1.000100E+4   1.311947E+0   7.329270E-5   
6.760950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.002000E+3   -9.002000E+3   1.186908E+0   7.189323E-5   
6.857550E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.001000E+3   -8.001000E+3   1.056461E+0   6.533169E-5   
6.954170E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.002000E+3   -7.002000E+3   9.217582E-1   5.426780E-5   
7.043090E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.002000E+3   -6.002000E+3   7.937722E-1   5.004428E-5   
7.139850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.001000E+3   -5.001000E+3   6.605758E-1   4.073403E-5   
7.231780E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.001000E+3   -4.001000E+3   5.298007E-1   3.372127E-5   
7.320730E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.002000E+3   -3.002000E+3   3.962100E-1   2.376915E-5   
7.412590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.001000E+3   -2.001000E+3   2.656530E-1   1.709835E-5   
7.504580E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.002000E+3   -1.002000E+3   1.298161E-1   4.899944E-6   
7.591140E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.000000E+0   -2.000000E+0   2.617691E-4   -8.919731E-7   
7.682030E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.960000E+2   9.960000E+2   -1.309068E-1   -8.545677E-6   
7.774490E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.998000E+3   1.998000E+3   -2.633843E-1   -1.701330E-5   
7.866860E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.997000E+3   2.997000E+3   -3.982823E-1   -2.827279E-5   
7.959290E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.998000E+3   3.998000E+3   -5.318295E-1   -3.793392E-5   
8.056660E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.998000E+3   4.998000E+3   -6.597045E-1   -4.204641E-5   
8.153990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.998000E+3   5.998000E+3   -7.862465E-1   -4.482589E-5   
8.251330E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.998000E+3   6.998000E+3   -9.171345E-1   -5.195154E-5   
8.343200E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.999000E+3   7.999000E+3   -1.055566E+0   -6.649689E-5   
8.440510E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.998000E+3   8.998000E+3   -1.171420E+0   -5.871210E-5   
8.532380E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.998000E+3   9.998000E+3   -1.312121E+0   -7.565093E-5   
8.627710E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.099800E+4   1.099800E+4   -1.443616E+0   -8.338325E-5   
8.726350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.199900E+4   1.199900E+4   -1.572123E+0   -8.800417E-5   
8.824990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.299800E+4   1.299800E+4   -1.699580E+0   -9.182209E-5   
8.923640E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.399800E+4   1.399800E+4   -1.823908E+0   -9.238806E-5   
9.027320E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499800E+4   1.499800E+4   -1.951977E+0   -9.669620E-5   
9.132910E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.599900E+4   1.599900E+4   -2.068005E+0   -9.122551E-5   
9.246550E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.699800E+4   1.699800E+4   -2.196467E+0   -1.005955E-4   
9.360250E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.799700E+4   1.799700E+4   -2.309749E+0   -9.702289E-5   
9.483960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.899700E+4   1.899700E+4   -2.428571E+0   -1.021295E-4   
@@END Data.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -364.655       -18997.000     9316.173       Coercive Field: Field at which M//H changes sign
Mr emu                                  -227.236E-9    907.311E-9     567.274E-9     Remanent Magnetization: M at H=0        
S                                       0.002          0.008          0.005          Squareness: Mr/Ms                       
S*                                      1.298          1.002          1.150          1-(Mr/Hc)(1/slope at Hc)                
M at H max emu                          -102.130E-6    96.662E-6      99.396E-6      M at the maximum field                  
                                                                                                                             

@END Measurement parameters
