@Filename: C:\vsm-lv\System_Admin\data\Dominique\DD146\empty_pot\empty_pot-Hys-00.VHD
@Measurement Controlfilename: c:\vsm-lv\System_Admin\Recipes\VC_HL_quickscan_allrange.VHC
@Calibration filename: c:\vsm-lv\System_Admin\settings\default.cal
@Parameter Filec:\vsm-lv\System_Admin\settings\default.cal
@Operator: System_Admin
@Samplename: empty_pot
@Date: Friday, September 30, 2016    (2016-09-30)
@Time: 14:44:28
@Test ID: test
@Apparatus: EZ7; LabVSM; Customer: Grubenhagen; first started on: Wednesday February 03, , 2015
[Installed Options]
VSM Model="EV X"
VSM=TRUE    
Torque=FALSE    
Signal Processor="SRS SR 830"
Torque Signal Processor="NI-6210"
Unipolar=FALSE    
Automation=FALSE    
MR=FALSE    
Torque Signal Inversion=TRUE    
VSM DAQ Card=TRUE    
Time Constant="0.1 s"
DAQ Output=FALSE    

[Signal and Coils]
Signal Connection="A-B"
Vector Coils=FALSE    
Stationary Coils=FALSE    
Z Coils=FALSE    
Sensor Angle="0 deg"
Time Between Averages=0.150000    
Y Averages Multiplier=1    
Reference Source="External"
SR830 Frequency=75.000000    

[Rotation]
Automatic Rotation=TRUE    
Rotate Option="Mdrive"
Rotation Display=FALSE    
Max Angle=400.000000    
Min Angle=-400.000000    
Rotation Serial Port=1    
Rotation Display Serial Port=1    
Torque Rotation Serial Port=4    

[Field]
Gaussmeter="32 KP DRC"
Gauss Probe="1 x"
Maximum Field=19000.000000    
Wait Time=4.000000    
Sweeprate Array="1500.000, 500.000, 100.000, 10.000, "
Averaging Array="1, 1, 1, 10, "
Precision Array="3.000, 0.500, 0.200, 0.200, "
Stability Array="1.000, 1.000, 0.500, 0.100, "
FCM-10 Address="GPIB0::16::INSTR"
Minimum Sweep Time=2.000000    
Minimum Sweep Rate Divider=40.000000    
Stability Time Between Readings=0.300000    
Number of Readings for Stability Check=2.000000    
Slow Approach=TRUE    
Slow Start %=90.000000    
Slow Approach Max Sweep Rate Divider=10.000000    
Max Slow Sweep Time=4.000000    

[MR]
MR Signal Processor=Manual VSM
Punch Through="Variable 0-10V"
Automation Comm Port=0
Max Current=20.000000    
Min AD Voltage=4.600000    
Max AD Voltage=7.000000    
MR Option=FALSE    
MS MR Signal Processor=FALSE    
AC&DC Current Source=FALSE    

[Temperature Control]
Temperature Control=TRUE    
Boil Off Nitrogen=FALSE    
Liquid Helium=FALSE    
Leave Temperature On=TRUE    
Temperature Control Type="SI 9700"
Sensor A="E-type"
Sensor B="E-type"
Control Sensor="A"
Sensor A Table=""
Sensor B Table=""
ITC Serial Port=2    
TC GPIB Address=15    
Temperature Log File="/c/vsm-lv/temperature.log"
Default Temperature=298.150000    
Gas Switching Temperature=333.150000    
Default Soak Time=120.000000    
Set Temperature Sample Time=10.000000    
Temperature Accuracy=1.000000    
Temperature Accuracy %=1.000000    
Automatic Gas Switching=FALSE    
1000 C Option=FALSE    
Number of points for accuracy wait=90    
Time between points for accuracy wait=1.000000    
Wait for Heat Exchanger Removal=FALSE    
Removal Temperature=0.000000    
Wait Time for Heat Exchanger Removal=0.000000    

[SI 9700]
P=1    
I=20    
D=0    
HE-P=1    
HE-I=20    
HE-D=0    
Max T Sweep Seed=1.000000
Min T Sweep Seed=0.200000
Max Heater Power=80    
Max T Sweep Speed=60.000000    
Min T Sweep Speed=12.000000    

[Other]
Transverse Direction="Absolute"
Default Transverse Direction=90.000000    
Time Dependence Start Field Distance=10.000000    
Minimum Remanence Wait Time=2.000000    
Default AC Demag Max Field=10000.000000    
AC Demag Minimum Field=1.000000    
Max Lockin Phase Error=90    
Mains Frequency=50.000000    
Samples Per Cycle=100    

[Interlock]
Door Lock=FALSE    
Interlock=FALSE    
Light Tower=FALSE    
Interlock Interface Name="Dev3"

[Torque Interface]
Torque Interface Name="Dev2"

[Exit Gas Heater Settings]
EGH PC Control=FALSE    
EGH Serial Port=0    
EGH Voltages=""

[VSM Interface]
VSM Interface Name="Dev1"

[MR Interface]
MR Interface Name="Dev1"

[DAQ Communication]
Protocol="Mx"
Remove Spikes=TRUE    

[Sensor Table]
1st Column=0    
Temperature Unit=0    

[Communication]
LIA 1 Address="GPIB0::8::INSTR"
LIA 2 Address=""
VSM Rotation Address="COM1"
Torque Rotation Address=""
Rotation Display Address=""
SI9700 Address="COM12"
EGH Address=""
Communication Mode="Original"
LIA Baud Rate="19200"
LIA Serial Read Delay=50    

[LIA]
Local=0    
Minimum Sensitivity="5 uV"

[MR External Current Source]
Ext I Src Adddress=""
AC MR Channel=""
DC MR Channel=""
Read Termination Character="CR"
CS Baud Rate="300"
Flow Control="Off"
Which LIA="1"
Input="A"
Ref Slope="Sine"
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Cylindrical;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 3.318E-7 [m^3] Area = 0.000E+0 [mm^2] Mass = 6.740E-3 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: MicroSense EasyVSM Software version EasyVSM 20150305-01
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to -0.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set VSM DAQ AO0 Voltage to 10.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 2:      Set VSM DAQ AO1 Voltage to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Applied Field to 0.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 4:      Set Auto Range Signal to 10.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = No
@Number of sections= 3
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From:  0.0000 [Oe] To: 19000.0000 [Oe] Min Stepsize/Sweeprate = 1000.0000 [Oe] Max Stepsize/Sweeprate = 1000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Measured Signal(s) = X
@Section 0 END
@Section 1: Hysteresis
@Preparation Actions: None
@Main Parameter Setup:
     From: 19000.0000 [Oe] To: -19000.0000 [Oe] Min Stepsize/Sweeprate = 1000.0000 [Oe] Max Stepsize/Sweeprate = 1000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: -19000.0000 [Oe] To: 19000.0000 [Oe] Min Stepsize/Sweeprate = 1000.0000 [Oe] Max Stepsize/Sweeprate = 1000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 2 END
@@Plot Settings
Number of plots: 1
Plot 0: Hysteresis = On; Section: 0; Signal: X; Label: Hys X; Point style: 2; Interpolation: On; Color: 14417948; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = FALSE
Sensor Angle = 0 deg
@Gauss Range: 30 kOe
@Emu Range: 5 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 5
@Rot 0 deg cal: -21170
@Rot 360 deg cal: 20810
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 10530
@Emu/v: 58.907
@Y Coils Correction Factor: 1.385
@Sample Shape Correction Factor: 1.000
@Coil Angle Alpha: 45.000
@Coil Angle Beta: -45.000
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 17
14998.000000   1.000000
15247.000000   1.000156
15497.000000   1.000302
15747.000000   1.000527
15997.000000   1.000751
16247.000000   1.001191
16497.000000   1.001494
16746.000000   1.001865
16996.000000   1.002237
17247.000000   1.002688
17496.000000   1.003286
17746.000000   1.003738
17996.000000   1.004259
18245.000000   1.005007
18495.000000   1.005686
18745.000000   1.006367
18995.000000   1.007118
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 0.700000
Background Subtraction = Yes   Method = Point by point
Background Signal array length = 32
-18993.000000   2.406274E-3   0.000000E+0   0.000000E+0
-18502.000000   2.348410E-3   0.000000E+0   0.000000E+0
-18001.000000   2.288960E-3   0.000000E+0   0.000000E+0
-17501.000000   2.227346E-3   0.000000E+0   0.000000E+0
-17002.000000   2.166318E-3   0.000000E+0   0.000000E+0
-16501.000000   2.104911E-3   0.000000E+0   0.000000E+0
-16000.000000   2.042623E-3   0.000000E+0   0.000000E+0
-15501.000000   1.978574E-3   0.000000E+0   0.000000E+0
-15001.000000   1.918608E-3   0.000000E+0   0.000000E+0
-13001.000000   1.670876E-3   0.000000E+0   0.000000E+0
-11001.000000   1.415849E-3   0.000000E+0   0.000000E+0
-9001.000000   1.161825E-3   0.000000E+0   0.000000E+0
-7002.000000   9.030077E-4   0.000000E+0   0.000000E+0
-5001.000000   6.471822E-4   0.000000E+0   0.000000E+0
-3002.000000   3.860235E-4   0.000000E+0   0.000000E+0
-1002.000000   1.238858E-4   0.000000E+0   0.000000E+0
995.000000   -1.233702E-4   0.000000E+0   0.000000E+0
2996.000000   -3.852079E-4   0.000000E+0   0.000000E+0
4997.000000   -6.443583E-4   0.000000E+0   0.000000E+0
6997.000000   -9.021850E-4   0.000000E+0   0.000000E+0
8998.000000   -1.158138E-3   0.000000E+0   0.000000E+0
10996.000000   -1.413947E-3   0.000000E+0   0.000000E+0
12997.000000   -1.666259E-3   0.000000E+0   0.000000E+0
14997.000000   -1.916258E-3   0.000000E+0   0.000000E+0
15498.000000   -1.978401E-3   0.000000E+0   0.000000E+0
15998.000000   -2.040843E-3   0.000000E+0   0.000000E+0
16498.000000   -2.100129E-3   0.000000E+0   0.000000E+0
16997.000000   -2.163433E-3   0.000000E+0   0.000000E+0
17498.000000   -2.225328E-3   0.000000E+0   0.000000E+0
17997.000000   -2.283674E-3   0.000000E+0   0.000000E+0
18496.000000   -2.348147E-3   0.000000E+0   0.000000E+0
18992.000000   -2.401551E-3   0.000000E+0   0.000000E+0
Angular Sensitivity Correction = Yes
Angular Sensitivity array length = 361
0.000000   1.000026E+0   0.000000E+0   0.000000
1.000000   9.998824E-1   0.000000E+0   0.000000
2.000000   9.997501E-1   0.000000E+0   0.000000
3.000000   9.996408E-1   0.000000E+0   0.000000
4.000000   9.995661E-1   0.000000E+0   0.000000
5.000000   9.995373E-1   0.000000E+0   0.000000
6.000000   9.995662E-1   0.000000E+0   0.000000
7.000000   9.996640E-1   0.000000E+0   0.000000
8.000000   9.998424E-1   0.000000E+0   0.000000
9.000000   1.000113E+0   0.000000E+0   0.000000
10.000000   1.000487E+0   0.000000E+0   0.000000
11.000000   1.000976E+0   0.000000E+0   0.000000
12.000000   1.001591E+0   0.000000E+0   0.000000
13.000000   1.002345E+0   0.000000E+0   0.000000
14.000000   1.003248E+0   0.000000E+0   0.000000
15.000000   1.004313E+0   0.000000E+0   0.000000
16.000000   1.005547E+0   0.000000E+0   0.000000
17.000000   1.006952E+0   0.000000E+0   0.000000
18.000000   1.008524E+0   0.000000E+0   0.000000
19.000000   1.010260E+0   0.000000E+0   0.000000
20.000000   1.012158E+0   0.000000E+0   0.000000
21.000000   1.014215E+0   0.000000E+0   0.000000
22.000000   1.016429E+0   0.000000E+0   0.000000
23.000000   1.018797E+0   0.000000E+0   0.000000
24.000000   1.021316E+0   0.000000E+0   0.000000
25.000000   1.023983E+0   0.000000E+0   0.000000
26.000000   1.026796E+0   0.000000E+0   0.000000
27.000000   1.029751E+0   0.000000E+0   0.000000
28.000000   1.032848E+0   0.000000E+0   0.000000
29.000000   1.036082E+0   0.000000E+0   0.000000
30.000000   1.039451E+0   0.000000E+0   0.000000
31.000000   1.042951E+0   0.000000E+0   0.000000
32.000000   1.046574E+0   0.000000E+0   0.000000
33.000000   1.050309E+0   0.000000E+0   0.000000
34.000000   1.054148E+0   0.000000E+0   0.000000
35.000000   1.058079E+0   0.000000E+0   0.000000
36.000000   1.062094E+0   0.000000E+0   0.000000
37.000000   1.066183E+0   0.000000E+0   0.000000
38.000000   1.070335E+0   0.000000E+0   0.000000
39.000000   1.074542E+0   0.000000E+0   0.000000
40.000000   1.078793E+0   0.000000E+0   0.000000
41.000000   1.083078E+0   0.000000E+0   0.000000
42.000000   1.087388E+0   0.000000E+0   0.000000
43.000000   1.091713E+0   0.000000E+0   0.000000
44.000000   1.096043E+0   0.000000E+0   0.000000
45.000000   1.100369E+0   0.000000E+0   0.000000
46.000000   1.104681E+0   0.000000E+0   0.000000
47.000000   1.108977E+0   0.000000E+0   0.000000
48.000000   1.113255E+0   0.000000E+0   0.000000
49.000000   1.117512E+0   0.000000E+0   0.000000
50.000000   1.121748E+0   0.000000E+0   0.000000
51.000000   1.125960E+0   0.000000E+0   0.000000
52.000000   1.130146E+0   0.000000E+0   0.000000
53.000000   1.134304E+0   0.000000E+0   0.000000
54.000000   1.138432E+0   0.000000E+0   0.000000
55.000000   1.142529E+0   0.000000E+0   0.000000
56.000000   1.146593E+0   0.000000E+0   0.000000
57.000000   1.150621E+0   0.000000E+0   0.000000
58.000000   1.154612E+0   0.000000E+0   0.000000
59.000000   1.158564E+0   0.000000E+0   0.000000
60.000000   1.162475E+0   0.000000E+0   0.000000
61.000000   1.166339E+0   0.000000E+0   0.000000
62.000000   1.170133E+0   0.000000E+0   0.000000
63.000000   1.173831E+0   0.000000E+0   0.000000
64.000000   1.177406E+0   0.000000E+0   0.000000
65.000000   1.180831E+0   0.000000E+0   0.000000
66.000000   1.184079E+0   0.000000E+0   0.000000
67.000000   1.187125E+0   0.000000E+0   0.000000
68.000000   1.189940E+0   0.000000E+0   0.000000
69.000000   1.192499E+0   0.000000E+0   0.000000
70.000000   1.194775E+0   0.000000E+0   0.000000
71.000000   1.196740E+0   0.000000E+0   0.000000
72.000000   1.198369E+0   0.000000E+0   0.000000
73.000000   1.199634E+0   0.000000E+0   0.000000
74.000000   1.200509E+0   0.000000E+0   0.000000
75.000000   1.200967E+0   0.000000E+0   0.000000
76.000000   1.200994E+0   0.000000E+0   0.000000
77.000000   1.200624E+0   0.000000E+0   0.000000
78.000000   1.199905E+0   0.000000E+0   0.000000
79.000000   1.198883E+0   0.000000E+0   0.000000
80.000000   1.197605E+0   0.000000E+0   0.000000
81.000000   1.196119E+0   0.000000E+0   0.000000
82.000000   1.194472E+0   0.000000E+0   0.000000
83.000000   1.192710E+0   0.000000E+0   0.000000
84.000000   1.190880E+0   0.000000E+0   0.000000
85.000000   1.189031E+0   0.000000E+0   0.000000
86.000000   1.187207E+0   0.000000E+0   0.000000
87.000000   1.185457E+0   0.000000E+0   0.000000
88.000000   1.183828E+0   0.000000E+0   0.000000
89.000000   1.182367E+0   0.000000E+0   0.000000
90.000000   1.181120E+0   0.000000E+0   0.000000
91.000000   1.180125E+0   0.000000E+0   0.000000
92.000000   1.179386E+0   0.000000E+0   0.000000
93.000000   1.178896E+0   0.000000E+0   0.000000
94.000000   1.178648E+0   0.000000E+0   0.000000
95.000000   1.178636E+0   0.000000E+0   0.000000
96.000000   1.178854E+0   0.000000E+0   0.000000
97.000000   1.179294E+0   0.000000E+0   0.000000
98.000000   1.179952E+0   0.000000E+0   0.000000
99.000000   1.180819E+0   0.000000E+0   0.000000
100.000000   1.181891E+0   0.000000E+0   0.000000
101.000000   1.183160E+0   0.000000E+0   0.000000
102.000000   1.184620E+0   0.000000E+0   0.000000
103.000000   1.186264E+0   0.000000E+0   0.000000
104.000000   1.188087E+0   0.000000E+0   0.000000
105.000000   1.190081E+0   0.000000E+0   0.000000
106.000000   1.192236E+0   0.000000E+0   0.000000
107.000000   1.194518E+0   0.000000E+0   0.000000
108.000000   1.196891E+0   0.000000E+0   0.000000
109.000000   1.199318E+0   0.000000E+0   0.000000
110.000000   1.201761E+0   0.000000E+0   0.000000
111.000000   1.204182E+0   0.000000E+0   0.000000
112.000000   1.206545E+0   0.000000E+0   0.000000
113.000000   1.208812E+0   0.000000E+0   0.000000
114.000000   1.210946E+0   0.000000E+0   0.000000
115.000000   1.212909E+0   0.000000E+0   0.000000
116.000000   1.214664E+0   0.000000E+0   0.000000
117.000000   1.216174E+0   0.000000E+0   0.000000
118.000000   1.217402E+0   0.000000E+0   0.000000
119.000000   1.218310E+0   0.000000E+0   0.000000
120.000000   1.218860E+0   0.000000E+0   0.000000
121.000000   1.219027E+0   0.000000E+0   0.000000
122.000000   1.218821E+0   0.000000E+0   0.000000
123.000000   1.218265E+0   0.000000E+0   0.000000
124.000000   1.217382E+0   0.000000E+0   0.000000
125.000000   1.216194E+0   0.000000E+0   0.000000
126.000000   1.214723E+0   0.000000E+0   0.000000
127.000000   1.212992E+0   0.000000E+0   0.000000
128.000000   1.211022E+0   0.000000E+0   0.000000
129.000000   1.208837E+0   0.000000E+0   0.000000
130.000000   1.206459E+0   0.000000E+0   0.000000
131.000000   1.203910E+0   0.000000E+0   0.000000
132.000000   1.201212E+0   0.000000E+0   0.000000
133.000000   1.198388E+0   0.000000E+0   0.000000
134.000000   1.195459E+0   0.000000E+0   0.000000
135.000000   1.192449E+0   0.000000E+0   0.000000
136.000000   1.189376E+0   0.000000E+0   0.000000
137.000000   1.186243E+0   0.000000E+0   0.000000
138.000000   1.183050E+0   0.000000E+0   0.000000
139.000000   1.179797E+0   0.000000E+0   0.000000
140.000000   1.176482E+0   0.000000E+0   0.000000
141.000000   1.173105E+0   0.000000E+0   0.000000
142.000000   1.169667E+0   0.000000E+0   0.000000
143.000000   1.166166E+0   0.000000E+0   0.000000
144.000000   1.162602E+0   0.000000E+0   0.000000
145.000000   1.158975E+0   0.000000E+0   0.000000
146.000000   1.155283E+0   0.000000E+0   0.000000
147.000000   1.151528E+0   0.000000E+0   0.000000
148.000000   1.147707E+0   0.000000E+0   0.000000
149.000000   1.143822E+0   0.000000E+0   0.000000
150.000000   1.139870E+0   0.000000E+0   0.000000
151.000000   1.135854E+0   0.000000E+0   0.000000
152.000000   1.131784E+0   0.000000E+0   0.000000
153.000000   1.127671E+0   0.000000E+0   0.000000
154.000000   1.123527E+0   0.000000E+0   0.000000
155.000000   1.119362E+0   0.000000E+0   0.000000
156.000000   1.115190E+0   0.000000E+0   0.000000
157.000000   1.111022E+0   0.000000E+0   0.000000
158.000000   1.106868E+0   0.000000E+0   0.000000
159.000000   1.102742E+0   0.000000E+0   0.000000
160.000000   1.098653E+0   0.000000E+0   0.000000
161.000000   1.094615E+0   0.000000E+0   0.000000
162.000000   1.090639E+0   0.000000E+0   0.000000
163.000000   1.086736E+0   0.000000E+0   0.000000
164.000000   1.082918E+0   0.000000E+0   0.000000
165.000000   1.079196E+0   0.000000E+0   0.000000
166.000000   1.075581E+0   0.000000E+0   0.000000
167.000000   1.072078E+0   0.000000E+0   0.000000
168.000000   1.068691E+0   0.000000E+0   0.000000
169.000000   1.065422E+0   0.000000E+0   0.000000
170.000000   1.062276E+0   0.000000E+0   0.000000
171.000000   1.059256E+0   0.000000E+0   0.000000
172.000000   1.056366E+0   0.000000E+0   0.000000
173.000000   1.053609E+0   0.000000E+0   0.000000
174.000000   1.050989E+0   0.000000E+0   0.000000
175.000000   1.048510E+0   0.000000E+0   0.000000
176.000000   1.046174E+0   0.000000E+0   0.000000
177.000000   1.043987E+0   0.000000E+0   0.000000
178.000000   1.041950E+0   0.000000E+0   0.000000
179.000000   1.040068E+0   0.000000E+0   0.000000
180.000000   1.038345E+0   0.000000E+0   0.000000
181.000000   1.036783E+0   0.000000E+0   0.000000
182.000000   1.035385E+0   0.000000E+0   0.000000
183.000000   1.034152E+0   0.000000E+0   0.000000
184.000000   1.033086E+0   0.000000E+0   0.000000
185.000000   1.032187E+0   0.000000E+0   0.000000
186.000000   1.031459E+0   0.000000E+0   0.000000
187.000000   1.030901E+0   0.000000E+0   0.000000
188.000000   1.030516E+0   0.000000E+0   0.000000
189.000000   1.030306E+0   0.000000E+0   0.000000
190.000000   1.030271E+0   0.000000E+0   0.000000
191.000000   1.030414E+0   0.000000E+0   0.000000
192.000000   1.030736E+0   0.000000E+0   0.000000
193.000000   1.031238E+0   0.000000E+0   0.000000
194.000000   1.031922E+0   0.000000E+0   0.000000
195.000000   1.032790E+0   0.000000E+0   0.000000
196.000000   1.033841E+0   0.000000E+0   0.000000
197.000000   1.035069E+0   0.000000E+0   0.000000
198.000000   1.036465E+0   0.000000E+0   0.000000
199.000000   1.038023E+0   0.000000E+0   0.000000
200.000000   1.039733E+0   0.000000E+0   0.000000
201.000000   1.041588E+0   0.000000E+0   0.000000
202.000000   1.043579E+0   0.000000E+0   0.000000
203.000000   1.045699E+0   0.000000E+0   0.000000
204.000000   1.047938E+0   0.000000E+0   0.000000
205.000000   1.050290E+0   0.000000E+0   0.000000
206.000000   1.052746E+0   0.000000E+0   0.000000
207.000000   1.055298E+0   0.000000E+0   0.000000
208.000000   1.057938E+0   0.000000E+0   0.000000
209.000000   1.060657E+0   0.000000E+0   0.000000
210.000000   1.063448E+0   0.000000E+0   0.000000
211.000000   1.066303E+0   0.000000E+0   0.000000
212.000000   1.069213E+0   0.000000E+0   0.000000
213.000000   1.072170E+0   0.000000E+0   0.000000
214.000000   1.075167E+0   0.000000E+0   0.000000
215.000000   1.078196E+0   0.000000E+0   0.000000
216.000000   1.081247E+0   0.000000E+0   0.000000
217.000000   1.084314E+0   0.000000E+0   0.000000
218.000000   1.087389E+0   0.000000E+0   0.000000
219.000000   1.090463E+0   0.000000E+0   0.000000
220.000000   1.093528E+0   0.000000E+0   0.000000
221.000000   1.096576E+0   0.000000E+0   0.000000
222.000000   1.099599E+0   0.000000E+0   0.000000
223.000000   1.102590E+0   0.000000E+0   0.000000
224.000000   1.105540E+0   0.000000E+0   0.000000
225.000000   1.108441E+0   0.000000E+0   0.000000
226.000000   1.111288E+0   0.000000E+0   0.000000
227.000000   1.114083E+0   0.000000E+0   0.000000
228.000000   1.116834E+0   0.000000E+0   0.000000
229.000000   1.119546E+0   0.000000E+0   0.000000
230.000000   1.122224E+0   0.000000E+0   0.000000
231.000000   1.124876E+0   0.000000E+0   0.000000
232.000000   1.127507E+0   0.000000E+0   0.000000
233.000000   1.130123E+0   0.000000E+0   0.000000
234.000000   1.132730E+0   0.000000E+0   0.000000
235.000000   1.135334E+0   0.000000E+0   0.000000
236.000000   1.137940E+0   0.000000E+0   0.000000
237.000000   1.140556E+0   0.000000E+0   0.000000
238.000000   1.143186E+0   0.000000E+0   0.000000
239.000000   1.145838E+0   0.000000E+0   0.000000
240.000000   1.148516E+0   0.000000E+0   0.000000
241.000000   1.151221E+0   0.000000E+0   0.000000
242.000000   1.153928E+0   0.000000E+0   0.000000
243.000000   1.156608E+0   0.000000E+0   0.000000
244.000000   1.159229E+0   0.000000E+0   0.000000
245.000000   1.161761E+0   0.000000E+0   0.000000
246.000000   1.164173E+0   0.000000E+0   0.000000
247.000000   1.166436E+0   0.000000E+0   0.000000
248.000000   1.168519E+0   0.000000E+0   0.000000
249.000000   1.170391E+0   0.000000E+0   0.000000
250.000000   1.172022E+0   0.000000E+0   0.000000
251.000000   1.173381E+0   0.000000E+0   0.000000
252.000000   1.174439E+0   0.000000E+0   0.000000
253.000000   1.175164E+0   0.000000E+0   0.000000
254.000000   1.175526E+0   0.000000E+0   0.000000
255.000000   1.175494E+0   0.000000E+0   0.000000
256.000000   1.175054E+0   0.000000E+0   0.000000
257.000000   1.174243E+0   0.000000E+0   0.000000
258.000000   1.173118E+0   0.000000E+0   0.000000
259.000000   1.171731E+0   0.000000E+0   0.000000
260.000000   1.170138E+0   0.000000E+0   0.000000
261.000000   1.168393E+0   0.000000E+0   0.000000
262.000000   1.166549E+0   0.000000E+0   0.000000
263.000000   1.164661E+0   0.000000E+0   0.000000
264.000000   1.162784E+0   0.000000E+0   0.000000
265.000000   1.160972E+0   0.000000E+0   0.000000
266.000000   1.159278E+0   0.000000E+0   0.000000
267.000000   1.157758E+0   0.000000E+0   0.000000
268.000000   1.156464E+0   0.000000E+0   0.000000
269.000000   1.155453E+0   0.000000E+0   0.000000
270.000000   1.154778E+0   0.000000E+0   0.000000
271.000000   1.154479E+0   0.000000E+0   0.000000
272.000000   1.154546E+0   0.000000E+0   0.000000
273.000000   1.154954E+0   0.000000E+0   0.000000
274.000000   1.155676E+0   0.000000E+0   0.000000
275.000000   1.156690E+0   0.000000E+0   0.000000
276.000000   1.157968E+0   0.000000E+0   0.000000
277.000000   1.159488E+0   0.000000E+0   0.000000
278.000000   1.161223E+0   0.000000E+0   0.000000
279.000000   1.163148E+0   0.000000E+0   0.000000
280.000000   1.165240E+0   0.000000E+0   0.000000
281.000000   1.167472E+0   0.000000E+0   0.000000
282.000000   1.169820E+0   0.000000E+0   0.000000
283.000000   1.172260E+0   0.000000E+0   0.000000
284.000000   1.174765E+0   0.000000E+0   0.000000
285.000000   1.177311E+0   0.000000E+0   0.000000
286.000000   1.179873E+0   0.000000E+0   0.000000
287.000000   1.182423E+0   0.000000E+0   0.000000
288.000000   1.184933E+0   0.000000E+0   0.000000
289.000000   1.187376E+0   0.000000E+0   0.000000
290.000000   1.189723E+0   0.000000E+0   0.000000
291.000000   1.191947E+0   0.000000E+0   0.000000
292.000000   1.194019E+0   0.000000E+0   0.000000
293.000000   1.195912E+0   0.000000E+0   0.000000
294.000000   1.197597E+0   0.000000E+0   0.000000
295.000000   1.199047E+0   0.000000E+0   0.000000
296.000000   1.200234E+0   0.000000E+0   0.000000
297.000000   1.201130E+0   0.000000E+0   0.000000
298.000000   1.201706E+0   0.000000E+0   0.000000
299.000000   1.201936E+0   0.000000E+0   0.000000
300.000000   1.201791E+0   0.000000E+0   0.000000
301.000000   1.201251E+0   0.000000E+0   0.000000
302.000000   1.200329E+0   0.000000E+0   0.000000
303.000000   1.199047E+0   0.000000E+0   0.000000
304.000000   1.197426E+0   0.000000E+0   0.000000
305.000000   1.195488E+0   0.000000E+0   0.000000
306.000000   1.193253E+0   0.000000E+0   0.000000
307.000000   1.190744E+0   0.000000E+0   0.000000
308.000000   1.187980E+0   0.000000E+0   0.000000
309.000000   1.184985E+0   0.000000E+0   0.000000
310.000000   1.181778E+0   0.000000E+0   0.000000
311.000000   1.178381E+0   0.000000E+0   0.000000
312.000000   1.174816E+0   0.000000E+0   0.000000
313.000000   1.171104E+0   0.000000E+0   0.000000
314.000000   1.167266E+0   0.000000E+0   0.000000
315.000000   1.163324E+0   0.000000E+0   0.000000
316.000000   1.159296E+0   0.000000E+0   0.000000
317.000000   1.155191E+0   0.000000E+0   0.000000
318.000000   1.151016E+0   0.000000E+0   0.000000
319.000000   1.146778E+0   0.000000E+0   0.000000
320.000000   1.142484E+0   0.000000E+0   0.000000
321.000000   1.138139E+0   0.000000E+0   0.000000
322.000000   1.133751E+0   0.000000E+0   0.000000
323.000000   1.129325E+0   0.000000E+0   0.000000
324.000000   1.124870E+0   0.000000E+0   0.000000
325.000000   1.120390E+0   0.000000E+0   0.000000
326.000000   1.115894E+0   0.000000E+0   0.000000
327.000000   1.111387E+0   0.000000E+0   0.000000
328.000000   1.106877E+0   0.000000E+0   0.000000
329.000000   1.102369E+0   0.000000E+0   0.000000
330.000000   1.097870E+0   0.000000E+0   0.000000
331.000000   1.093388E+0   0.000000E+0   0.000000
332.000000   1.088932E+0   0.000000E+0   0.000000
333.000000   1.084513E+0   0.000000E+0   0.000000
334.000000   1.080140E+0   0.000000E+0   0.000000
335.000000   1.075824E+0   0.000000E+0   0.000000
336.000000   1.071575E+0   0.000000E+0   0.000000
337.000000   1.067403E+0   0.000000E+0   0.000000
338.000000   1.063319E+0   0.000000E+0   0.000000
339.000000   1.059332E+0   0.000000E+0   0.000000
340.000000   1.055454E+0   0.000000E+0   0.000000
341.000000   1.051693E+0   0.000000E+0   0.000000
342.000000   1.048060E+0   0.000000E+0   0.000000
343.000000   1.044566E+0   0.000000E+0   0.000000
344.000000   1.041221E+0   0.000000E+0   0.000000
345.000000   1.038035E+0   0.000000E+0   0.000000
346.000000   1.035014E+0   0.000000E+0   0.000000
347.000000   1.032151E+0   0.000000E+0   0.000000
348.000000   1.029434E+0   0.000000E+0   0.000000
349.000000   1.026853E+0   0.000000E+0   0.000000
350.000000   1.024396E+0   0.000000E+0   0.000000
351.000000   1.022052E+0   0.000000E+0   0.000000
352.000000   1.019809E+0   0.000000E+0   0.000000
353.000000   1.017656E+0   0.000000E+0   0.000000
354.000000   1.015583E+0   0.000000E+0   0.000000
355.000000   1.013576E+0   0.000000E+0   0.000000
356.000000   1.011627E+0   0.000000E+0   0.000000
357.000000   1.009722E+0   0.000000E+0   0.000000
358.000000   1.007851E+0   0.000000E+0   0.000000
359.000000   1.006003E+0   0.000000E+0   0.000000
360.000000   1.004166E+0   0.000000E+0   0.000000
Remove Slope = No

Remove Signal Offset = No
Remove Signal Drift = FALSE; Drift # Points = 0
Remove Field Offset = No
Field Offset Method = Automatic
Field Offset = 0.0000
Remove Field Lag = No
Field Lag Method = Automatic
Field Lag = 0.0000
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0   Filter Type = Median
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = Thursday, September 01, 2016  17:19:09
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 3
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Temperature 2, Sample Temperature [degC]
Column 4: Raw Applied Field, Applied Field [Oe]
Column 5: Applied Field, Applied Field [Oe]
Column 6: Field Angle, Field Angle [deg]
Column 7: Raw Applied Field For Plot , Applied Field [Oe]
Column 8: Applied Field For Plot , Applied Field [Oe]
Column 9: Raw Signal Mx, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Temperature_2   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Signal_X_direction      
@Time at start of measurement: 14:44:29
@@Data
New Section: Section 0: 
3.560000E+0   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   1.124676E-4   2.880186E-7   
1.285800E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.980000E+2   9.980000E+2   -1.244935E-1   -7.339377E-7   
2.185800E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.999000E+3   1.999000E+3   -2.508576E-1   3.882926E-6   
3.202400E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.999000E+3   2.999000E+3   -3.787408E-1   6.845761E-6   
4.072600E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.999000E+3   3.999000E+3   -5.063513E-1   8.742395E-6   
5.085400E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.999000E+3   4.999000E+3   -6.310030E-1   1.359672E-5   
6.003800E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.999000E+3   5.999000E+3   -7.600717E-1   1.343802E-5   
6.923300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.999000E+3   6.999000E+3   -8.879210E-1   1.449674E-5   
7.837800E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.000000E+3   8.000000E+3   -1.014249E+0   1.620560E-5   
8.747300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.000000E+3   9.000000E+3   -1.139336E+0   1.902859E-5   
9.751600E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000000E+4   1.000000E+4   -1.267688E+0   1.870542E-5   
1.067890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100000E+4   1.100000E+4   -1.394992E+0   1.942306E-5   
1.160480E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200000E+4   1.200000E+4   -1.514436E+0   2.606853E-5   
1.253360E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300000E+4   1.300000E+4   -1.642329E+0   2.426198E-5   
1.345980E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400000E+4   1.400000E+4   -1.764432E+0   2.715602E-5   
1.441370E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499900E+4   1.499900E+4   -1.881228E+0   3.522848E-5   
1.539140E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600000E+4   1.600000E+4   -2.006556E+0   3.295485E-5   
1.647020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700000E+4   1.700000E+4   -2.125385E+0   3.359353E-5   
1.760280E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.800000E+4   1.800000E+4   -2.243031E+0   3.139154E-5   
1.883090E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.900000E+4   1.900000E+4   -2.348717E+0   3.605390E-5   
2.009690E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.800700E+4   1.800700E+4   -2.241846E+0   3.343914E-5   
2.127960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700500E+4   1.700500E+4   -2.127053E+0   3.252008E-5   
2.236590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600600E+4   1.600600E+4   -2.004117E+0   3.608579E-5   
2.344670E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.500500E+4   1.500500E+4   -1.884278E+0   3.291531E-5   
2.443340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400600E+4   1.400600E+4   -1.759494E+0   3.284377E-5   
2.541590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300400E+4   1.300400E+4   -1.636688E+0   3.040311E-5   
2.640350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200500E+4   1.200500E+4   -1.521019E+0   2.011650E-5   
2.739270E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100400E+4   1.100400E+4   -1.394070E+0   2.084995E-5   
2.832830E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000500E+4   1.000500E+4   -1.266527E+0   2.050726E-5   
2.929930E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.004000E+3   9.004000E+3   -1.142846E+0   1.603092E-5   
3.026950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.004000E+3   8.004000E+3   -1.017565E+0   1.340185E-5   
3.123930E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.003000E+3   7.003000E+3   -8.891180E-1   1.381136E-5   
3.220970E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.003000E+3   6.003000E+3   -7.581713E-1   1.585408E-5   
3.317960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.002000E+3   5.002000E+3   -6.340744E-1   1.091194E-5   
3.410290E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.004000E+3   4.004000E+3   -5.093851E-1   6.356133E-6   
3.502450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.003000E+3   3.003000E+3   -3.814673E-1   4.637257E-6   
3.594650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.004000E+3   2.004000E+3   -2.497989E-1   5.595906E-6   
3.687020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.002000E+3   1.002000E+3   -1.217723E-1   2.510720E-6   
3.776540E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.000000E+0   3.000000E+0   -2.413935E-3   -1.867009E-6   
3.867620E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.960000E+2   -9.960000E+2   1.240545E-1   9.147901E-7   
3.959960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.995000E+3   -1.995000E+3   2.537270E-1   -3.035981E-7   
4.052450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.996000E+3   -2.996000E+3   3.735892E-1   -1.163813E-5   
4.144840E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.995000E+3   -3.995000E+3   5.053691E-1   -1.037143E-5   
4.242300E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.997000E+3   -4.997000E+3   6.422378E-1   -4.405083E-6   
4.339300E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.997000E+3   -5.997000E+3   7.613759E-1   -1.312393E-5   
4.436130E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.997000E+3   -6.997000E+3   8.849038E-1   -1.744170E-5   
4.533080E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.997000E+3   -7.997000E+3   1.013350E+0   -1.845699E-5   
4.629990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.997000E+3   -8.997000E+3   1.148968E+0   -1.230883E-5   
4.726950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.997000E+3   -9.997000E+3   1.260821E+0   -2.747539E-5   
4.822450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.099700E+4   -1.099700E+4   1.387070E+0   -2.823473E-5   
4.921260E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.199800E+4   -1.199800E+4   1.510508E+0   -3.243221E-5   
5.020040E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.299800E+4   -1.299800E+4   1.637480E+0   -3.297083E-5   
5.118850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.399600E+4   -1.399600E+4   1.764672E+0   -2.940484E-5   
5.217650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.499600E+4   -1.499600E+4   1.890401E+0   -2.753894E-5   
5.326220E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.599700E+4   -1.599700E+4   2.002494E+0   -3.818747E-5   
5.440230E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.699800E+4   -1.699800E+4   2.126087E+0   -3.492149E-5   
5.559170E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.799700E+4   -1.799700E+4   2.241605E+0   -3.725009E-5   
5.683030E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.899800E+4   -1.899800E+4   2.346523E+0   -4.298748E-5   
5.814750E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.800300E+4   -1.800300E+4   2.236316E+0   -4.325141E-5   
5.928190E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.700300E+4   -1.700300E+4   2.121018E+0   -4.059608E-5   
6.026680E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.600400E+4   -1.600400E+4   2.004579E+0   -3.695938E-5   
6.130000E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.500300E+4   -1.500300E+4   1.879231E+0   -3.956257E-5   
6.228420E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.400200E+4   -1.400200E+4   1.766429E+0   -2.839137E-5   
6.331850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.300200E+4   -1.300200E+4   1.635923E+0   -3.503479E-5   
6.427300E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.200100E+4   -1.200100E+4   1.519067E+0   -2.425645E-5   
6.525950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.100100E+4   -1.100100E+4   1.388232E+0   -2.758109E-5   
6.620950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000000E+4   -1.000000E+4   1.264002E+0   -2.467533E-5   
6.709860E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.001000E+3   -9.001000E+3   1.140849E+0   -2.094675E-5   
6.798660E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.001000E+3   -8.001000E+3   1.019188E+0   -1.313700E-5   
6.892290E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.001000E+3   -7.001000E+3   8.884818E-1   -1.437496E-5   
6.978750E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.001000E+3   -6.001000E+3   7.596876E-1   -1.532366E-5   
7.067770E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.001000E+3   -5.001000E+3   6.343372E-1   -1.282854E-5   
7.154000E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.000000E+3   -4.000000E+3   5.085291E-1   -7.864535E-6   
7.240330E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.001000E+3   -3.001000E+3   3.812041E-1   -4.678421E-6   
7.326360E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.000000E+3   -2.000000E+3   2.513789E-1   -3.307056E-6   
7.415390E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.001000E+3   -1.001000E+3   1.244496E-1   6.908833E-7   
7.498380E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000000E+0   -1.000000E+0   2.194422E-5   7.367909E-8   
7.590460E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.980000E+2   9.980000E+2   -1.192707E-1   4.488937E-6   
7.677440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.999000E+3   1.999000E+3   -2.534416E-1   1.298822E-6   
7.769810E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.999000E+3   2.999000E+3   -3.772539E-1   8.332743E-6   
7.856800E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.999000E+3   3.999000E+3   -5.140813E-1   1.012234E-6   
7.948690E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.999000E+3   4.999000E+3   -6.292464E-1   1.535339E-5   
8.040270E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.000000E+3   6.000000E+3   -7.623856E-1   1.125299E-5   
8.131710E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.999000E+3   6.999000E+3   -8.854092E-1   1.700863E-5   
8.223340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.001000E+3   8.001000E+3   -1.008961E+0   2.162237E-5   
8.314150E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.000000E+3   9.000000E+3   -1.133848E+0   2.451656E-5   
8.405460E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000000E+4   1.000000E+4   -1.258473E+0   2.792114E-5   
8.498030E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100000E+4   1.100000E+4   -1.394178E+0   2.023718E-5   
8.590660E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200000E+4   1.200000E+4   -1.516039E+0   2.446620E-5   
8.683520E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300000E+4   1.300000E+4   -1.640926E+0   2.566519E-5   
8.776120E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400000E+4   1.400000E+4   -1.765155E+0   2.643261E-5   
8.871630E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499900E+4   1.499900E+4   -1.878395E+0   3.806083E-5   
8.969440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600000E+4   1.600000E+4   -2.007608E+0   3.190194E-5   
9.077240E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700000E+4   1.700000E+4   -2.119460E+0   3.953189E-5   
9.190510E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.800000E+4   1.800000E+4   -2.239278E+0   3.516126E-5   
9.309260E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.899900E+4   1.899900E+4   -2.347159E+0   3.762373E-5   
@@END Data.
@Time at end of measurement: 15:00:03
@Instrument  Changes:
@Emu Range: 50 uV
@END Instrument  Changes:
First Error: 2016-09-30  09:44:05
32KP Set Field V2

Set Field: Field did not reach target field Target = 20000.000000, Reached = 19000.000000
Start Field18999.000 [Oe]   Field to set 20000.000 [Oe]   Limited Field 19000.000 [Oe]   
Timer at start = 2110169, Timer now = 2112308, difference = 2139, total sweep time + 100 = 767
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = 19000.000
 Timer Now = 2112308
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19000.000
19000.000
 Timer Now = 2112308

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19000.000
19000.000
 Timer Now = 2112308
Error History:
Actions History:
2016-09-30  09:44:05
32KP Set Field V2

Set Field: Field did not reach target field Target = 20000.000000, Reached = 19000.000000
Start Field18999.000 [Oe]   Field to set 20000.000 [Oe]   Limited Field 19000.000 [Oe]   
Timer at start = 2110169, Timer now = 2112308, difference = 2139, total sweep time + 100 = 767
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = 19000.000
 Timer Now = 2112308
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19000.000
19000.000
 Timer Now = 2112308

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19000.000
19000.000
 Timer Now = 2112308

2016-09-30  10:02:14
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -18999.000000
Start Field-18999.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 3199402, Timer now = 3201554, difference = 2152, total sweep time + 100 = 767
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -18999.000
 Timer Now = 3201554
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -18999.000
-18999.000
 Timer Now = 3201554

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -18999.000
-18999.000
 Timer Now = 3201554

2016-09-30  10:02:45
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -18999.000000
Start Field-19000.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 3230966, Timer now = 3233028, difference = 2062, total sweep time + 100 = 100
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -18999.000
 Timer Now = 3233028
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -18999.000
-18999.000
 Timer Now = 3233028

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -18999.000
-18999.000
 Timer Now = 3233028

2016-09-30  10:03:10
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -18999.000000
Start Field-18999.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 3254949, Timer now = 3257104, difference = 2155, total sweep time + 100 = 767
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -18999.000
 Timer Now = 3257104
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -18999.000
-18999.000
 Timer Now = 3257104

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -18999.000
-18999.000
 Timer Now = 3257104

2016-09-30  10:31:00
32KP Set Field V2

Set Field: Field did not reach target field Target = 20000.000000, Reached = 19002.000000
Start Field19001.000 [Oe]   Field to set 20000.000 [Oe]   Limited Field 19000.000 [Oe]   
Timer at start = 4925033, Timer now = 4927169, difference = 2136, total sweep time + 100 = 767
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = 19002.000
 Timer Now = 4927169
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19002.000
19002.000
 Timer Now = 4927169

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19002.000
19002.000
 Timer Now = 4927169

2016-09-30  10:49:21
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -19000.000000
Start Field-18999.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 6026443, Timer now = 6028583, difference = 2140, total sweep time + 100 = 767
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -19000.000
 Timer Now = 6028583
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 6028583

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 6028583

2016-09-30  10:49:51
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -19000.000000
Start Field-19000.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 6056803, Timer now = 6058863, difference = 2060, total sweep time + 100 = 100
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -19000.000
 Timer Now = 6058863
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 6058863

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 6058863

2016-09-30  10:50:15
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -19000.000000
Start Field-19000.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 6080458, Timer now = 6082534, difference = 2076, total sweep time + 100 = 100
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -19000.000
 Timer Now = 6082534
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 6082534

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 6082534

2016-09-30  11:07:29
32KP Set Field V2

Set Field: Field did not reach target field Target = 20000.000000, Reached = 19002.000000
Start Field19002.000 [Oe]   Field to set 20000.000 [Oe]   Limited Field 19000.000 [Oe]   
Timer at start = 7114734, Timer now = 7116886, difference = 2152, total sweep time + 100 = 773
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = 19002.000
 Timer Now = 7116886
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19002.000
19002.000
 Timer Now = 7116886

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19002.000
19002.000
 Timer Now = 7116886

2016-09-30  11:25:08
32KP Set Field V2

Set Field: Field did not reach target field Target = 20000.000000, Reached = 19002.000000
Start Field19002.000 [Oe]   Field to set 20000.000 [Oe]   Limited Field 19000.000 [Oe]   
Timer at start = 8173294, Timer now = 8175430, difference = 2136, total sweep time + 100 = 773
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = 19002.000
 Timer Now = 8175430
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19002.000
19002.000
 Timer Now = 8175430

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19002.000
19002.000
 Timer Now = 8175430

2016-09-30  11:43:35
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -19000.000000
Start Field-19000.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 9280854, Timer now = 9282914, difference = 2060, total sweep time + 100 = 100
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -19000.000
 Timer Now = 9282914
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 9282914

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 9282914

2016-09-30  11:44:02
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -19000.000000
Start Field-19001.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 9307477, Timer now = 9309619, difference = 2142, total sweep time + 100 = 767
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -19000.000
 Timer Now = 9309619
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 9309619

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 9309619

2016-09-30  11:44:25
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -19000.000000
Start Field-19000.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 9330458, Timer now = 9332519, difference = 2061, total sweep time + 100 = 100
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -19000.000
 Timer Now = 9332519
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 9332519

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 9332519

2016-09-30  12:01:41
32KP Set Field V2

Set Field: Field did not reach target field Target = 20000.000000, Reached = 19002.000000
Start Field19002.000 [Oe]   Field to set 20000.000 [Oe]   Limited Field 19000.000 [Oe]   
Timer at start = 10366049, Timer now = 10368185, difference = 2136, total sweep time + 100 = 773
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = 19002.000
 Timer Now = 10368185
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19002.000
19002.000
 Timer Now = 10368185

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19002.000
19002.000
 Timer Now = 10368185

2016-09-30  13:10:59
32KP Set Field V2

Set Field: Field did not reach target field Target = 20000.000000, Reached = 19003.000000
Start Field19002.000 [Oe]   Field to set 20000.000 [Oe]   Limited Field 19000.000 [Oe]   
Timer at start = 14524875, Timer now = 14527027, difference = 2152, total sweep time + 100 = 773
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = 19003.000
 Timer Now = 14527027
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19003.000
19003.000
 Timer Now = 14527027

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19003.000
19003.000
 Timer Now = 14527027

2016-09-30  13:29:28
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -19000.000000
Start Field-19000.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 15633446, Timer now = 15635516, difference = 2070, total sweep time + 100 = 100
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -19000.000
 Timer Now = 15635516
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 15635516

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19000.000
-19000.000
 Timer Now = 15635516

2016-09-30  13:29:57
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -19001.000000
Start Field-19000.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 15662727, Timer now = 15664789, difference = 2062, total sweep time + 100 = 100
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -19001.000
 Timer Now = 15664789
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19001.000
-19000.000
 Timer Now = 15664789

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19001.000
-19000.000
 Timer Now = 15664789

2016-09-30  13:30:20
32KP Set Field V2

Set Field: Field did not reach target field Target = -20000.000000, Reached = -19001.000000
Start Field-19001.000 [Oe]   Field to set -20000.000 [Oe]   Limited Field -19000.000 [Oe]   
Timer at start = 15685825, Timer now = 15687974, difference = 2149, total sweep time + 100 = 767
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = -19001.000
 Timer Now = 15687974
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19001.000
-19000.000
 Timer Now = 15687974

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = TRUE; Stable=  TRUE; Stability Array = -19001.000
-19000.000
 Timer Now = 15687974

2016-09-30  13:47:34
32KP Set Field V2

Set Field: Field did not reach target field Target = 20000.000000, Reached = 19003.000000
Start Field19003.000 [Oe]   Field to set 20000.000 [Oe]   Limited Field 19000.000 [Oe]   
Timer at start = 16719735, Timer now = 16721874, difference = 2139, total sweep time + 100 = 780
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  FALSE; Stability Array = 19003.000
 Timer Now = 16721874
Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19003.000
19002.000
 Timer Now = 16721874

Reason wait ended:Stop Global = FALSE; Decreased Precision = FALSE; Slow Approach = FALSE; >=20 seconds =  FALSE; Field reached = FALSE; Stable=  TRUE; Stability Array = 19003.000
19002.000
 Timer Now = 16721874

@@Final Manipulated Data
New Section: Section 0: 
3.560000E+0   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   1.124676E-4   2.880186E-7   
1.285800E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.980000E+2   9.980000E+2   -1.244935E-1   -7.339377E-7   
2.185800E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.999000E+3   1.999000E+3   -2.508576E-1   3.882926E-6   
3.202400E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.999000E+3   2.999000E+3   -3.787408E-1   6.845761E-6   
4.072600E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.999000E+3   3.999000E+3   -5.063513E-1   8.742395E-6   
5.085400E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.999000E+3   4.999000E+3   -6.310030E-1   1.359672E-5   
6.003800E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.999000E+3   5.999000E+3   -7.600717E-1   1.343802E-5   
6.923300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.999000E+3   6.999000E+3   -8.879210E-1   1.449674E-5   
7.837800E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.000000E+3   8.000000E+3   -1.014249E+0   1.620560E-5   
8.747300E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.000000E+3   9.000000E+3   -1.139336E+0   1.902859E-5   
9.751600E+1   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000000E+4   1.000000E+4   -1.267688E+0   1.870542E-5   
1.067890E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100000E+4   1.100000E+4   -1.394992E+0   1.942306E-5   
1.160480E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200000E+4   1.200000E+4   -1.514436E+0   2.606853E-5   
1.253360E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300000E+4   1.300000E+4   -1.642329E+0   2.426198E-5   
1.345980E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400000E+4   1.400000E+4   -1.764432E+0   2.715602E-5   
1.441370E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499900E+4   1.499900E+4   -1.881228E+0   3.522848E-5   
1.539140E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600000E+4   1.600000E+4   -2.006556E+0   3.295485E-5   
1.647020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700000E+4   1.700000E+4   -2.125385E+0   3.359353E-5   
1.760280E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.800000E+4   1.800000E+4   -2.243031E+0   3.139154E-5   
1.883090E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.900000E+4   1.900000E+4   -2.348717E+0   3.605390E-5   
2.009690E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.800700E+4   1.800700E+4   -2.241846E+0   3.343914E-5   
2.127960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700500E+4   1.700500E+4   -2.127053E+0   3.252008E-5   
2.236590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600600E+4   1.600600E+4   -2.004117E+0   3.608579E-5   
2.344670E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.500500E+4   1.500500E+4   -1.884278E+0   3.291531E-5   
2.443340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400600E+4   1.400600E+4   -1.759494E+0   3.284377E-5   
2.541590E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300400E+4   1.300400E+4   -1.636688E+0   3.040311E-5   
2.640350E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200500E+4   1.200500E+4   -1.521019E+0   2.011650E-5   
2.739270E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100400E+4   1.100400E+4   -1.394070E+0   2.084995E-5   
2.832830E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000500E+4   1.000500E+4   -1.266527E+0   2.050726E-5   
2.929930E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.004000E+3   9.004000E+3   -1.142846E+0   1.603092E-5   
3.026950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.004000E+3   8.004000E+3   -1.017565E+0   1.340185E-5   
3.123930E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   7.003000E+3   7.003000E+3   -8.891180E-1   1.381136E-5   
3.220970E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.003000E+3   6.003000E+3   -7.581713E-1   1.585408E-5   
3.317960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   5.002000E+3   5.002000E+3   -6.340744E-1   1.091194E-5   
3.410290E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.004000E+3   4.004000E+3   -5.093851E-1   6.356133E-6   
3.502450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.003000E+3   3.003000E+3   -3.814673E-1   4.637257E-6   
3.594650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.004000E+3   2.004000E+3   -2.497989E-1   5.595906E-6   
3.687020E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.002000E+3   1.002000E+3   -1.217723E-1   2.510720E-6   
3.776540E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.000000E+0   3.000000E+0   -2.413935E-3   -1.867009E-6   
3.867620E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.960000E+2   -9.960000E+2   1.240545E-1   9.147901E-7   
3.959960E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.995000E+3   -1.995000E+3   2.537270E-1   -3.035981E-7   
4.052450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.996000E+3   -2.996000E+3   3.735892E-1   -1.163813E-5   
4.144840E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.995000E+3   -3.995000E+3   5.053691E-1   -1.037143E-5   
4.242300E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.997000E+3   -4.997000E+3   6.422378E-1   -4.405083E-6   
4.339300E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.997000E+3   -5.997000E+3   7.613759E-1   -1.312393E-5   
4.436130E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.997000E+3   -6.997000E+3   8.849038E-1   -1.744170E-5   
4.533080E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.997000E+3   -7.997000E+3   1.013350E+0   -1.845699E-5   
4.629990E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.997000E+3   -8.997000E+3   1.148968E+0   -1.230883E-5   
4.726950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.997000E+3   -9.997000E+3   1.260821E+0   -2.747539E-5   
4.822450E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.099700E+4   -1.099700E+4   1.387070E+0   -2.823473E-5   
4.921260E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.199800E+4   -1.199800E+4   1.510508E+0   -3.243221E-5   
5.020040E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.299800E+4   -1.299800E+4   1.637480E+0   -3.297083E-5   
5.118850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.399600E+4   -1.399600E+4   1.764672E+0   -2.940484E-5   
5.217650E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.499600E+4   -1.499600E+4   1.890401E+0   -2.753894E-5   
5.326220E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.599700E+4   -1.599700E+4   2.002494E+0   -3.818747E-5   
5.440230E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.699800E+4   -1.699800E+4   2.126087E+0   -3.492149E-5   
5.559170E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.799700E+4   -1.799700E+4   2.241605E+0   -3.725009E-5   
5.683030E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.899800E+4   -1.899800E+4   2.346523E+0   -4.298748E-5   
5.814750E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.800300E+4   -1.800300E+4   2.236316E+0   -4.325141E-5   
5.928190E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.700300E+4   -1.700300E+4   2.121018E+0   -4.059608E-5   
6.026680E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.600400E+4   -1.600400E+4   2.004579E+0   -3.695938E-5   
6.130000E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.500300E+4   -1.500300E+4   1.879231E+0   -3.956257E-5   
6.228420E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.400200E+4   -1.400200E+4   1.766429E+0   -2.839137E-5   
6.331850E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.300200E+4   -1.300200E+4   1.635923E+0   -3.503479E-5   
6.427300E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.200100E+4   -1.200100E+4   1.519067E+0   -2.425645E-5   
6.525950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.100100E+4   -1.100100E+4   1.388232E+0   -2.758109E-5   
6.620950E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000000E+4   -1.000000E+4   1.264002E+0   -2.467533E-5   
6.709860E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -9.001000E+3   -9.001000E+3   1.140849E+0   -2.094675E-5   
6.798660E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -8.001000E+3   -8.001000E+3   1.019188E+0   -1.313700E-5   
6.892290E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -7.001000E+3   -7.001000E+3   8.884818E-1   -1.437496E-5   
6.978750E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -6.001000E+3   -6.001000E+3   7.596876E-1   -1.532366E-5   
7.067770E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -5.001000E+3   -5.001000E+3   6.343372E-1   -1.282854E-5   
7.154000E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -4.000000E+3   -4.000000E+3   5.085291E-1   -7.864535E-6   
7.240330E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -3.001000E+3   -3.001000E+3   3.812041E-1   -4.678421E-6   
7.326360E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -2.000000E+3   -2.000000E+3   2.513789E-1   -3.307056E-6   
7.415390E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.001000E+3   -1.001000E+3   1.244496E-1   6.908833E-7   
7.498380E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   -1.000000E+0   -1.000000E+0   2.194422E-5   7.367909E-8   
7.590460E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.980000E+2   9.980000E+2   -1.192707E-1   4.488937E-6   
7.677440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.999000E+3   1.999000E+3   -2.534416E-1   1.298822E-6   
7.769810E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   2.999000E+3   2.999000E+3   -3.772539E-1   8.332743E-6   
7.856800E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   3.999000E+3   3.999000E+3   -5.140813E-1   1.012234E-6   
7.948690E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   4.999000E+3   4.999000E+3   -6.292464E-1   1.535339E-5   
8.040270E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.000000E+3   6.000000E+3   -7.623856E-1   1.125299E-5   
8.131710E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   6.999000E+3   6.999000E+3   -8.854092E-1   1.700863E-5   
8.223340E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   8.001000E+3   8.001000E+3   -1.008961E+0   2.162237E-5   
8.314150E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   9.000000E+3   9.000000E+3   -1.133848E+0   2.451656E-5   
8.405460E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.000000E+4   1.000000E+4   -1.258473E+0   2.792114E-5   
8.498030E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.100000E+4   1.100000E+4   -1.394178E+0   2.023718E-5   
8.590660E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.200000E+4   1.200000E+4   -1.516039E+0   2.446620E-5   
8.683520E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.300000E+4   1.300000E+4   -1.640926E+0   2.566519E-5   
8.776120E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.400000E+4   1.400000E+4   -1.765155E+0   2.643261E-5   
8.871630E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.499900E+4   1.499900E+4   -1.878395E+0   3.806083E-5   
8.969440E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.600000E+4   1.600000E+4   -2.007608E+0   3.190194E-5   
9.077240E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.700000E+4   1.700000E+4   -2.119460E+0   3.953189E-5   
9.190510E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.800000E+4   1.800000E+4   -2.239278E+0   3.516126E-5   
9.309260E+2   -2.731500E+2   -2.731500E+2   -2.731500E+2   0.000000E+0   0.000000E+0   0.000000E+0   1.899900E+4   1.899900E+4   -2.347159E+0   3.762373E-5   
@@END Data.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -281.267       18999.000      -9640.133      Coercive Field: Field at which M//H changes sign
Mr emu                                  -288.019E-9    37.624E-6      18.956E-6      Remanent Magnetization: M at H=0        
S                                       0.007          0.870          0.439          Squareness: Mr/Ms                       
S*                                      46.859         0.997          23.928         1-(Mr/Hc)(1/slope at Hc)                
M at H max emu                          36.054E-6      -42.987E-6     39.521E-6      M at the maximum field                  
                                                                                                                             

@END Measurement parameters
